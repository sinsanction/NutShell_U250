//commit c9a33ad89d777d8483ea4a2af9771f8176ba29bb
//Author: sinsanction <1602723930@qq.com>
//Date:   Mon Sep 12 10:29:22 2022 +0800
//
//    test cnnapibench lenet5 real func
//diff --git a/Makefile b/Makefile
//index 69ad24a..add34af 100644
//--- a/Makefile
//+++ b/Makefile
//@@ -11,7 +11,7 @@ SIMTOP = top.TopMain
// IMAGE ?= ready-to-run/linux.bin
// 
// DATAWIDTH ?= 64
//-BOARD ?= sim  # sim  pynq  axu3cg
//+BOARD ?= pynq  # sim  pynq  axu3cg
// CORE  ?= inorder  # inorder  ooo  embedded
// 
// .DEFAULT_GOAL = verilog
//diff --git a/src/main/scala/top/Settings.scala b/src/main/scala/top/Settings.scala
//index 9464530..18ee3af 100644
//--- a/src/main/scala/top/Settings.scala
//+++ b/src/main/scala/top/Settings.scala
//@@ -48,11 +48,11 @@ object PynqSettings {
//   def apply() = Map(
//     "FPGAPlatform" -> true,
//     "NrExtIntr" -> 3,
//-    "ResetVector" -> 0x60000000L,
//-    "MemMapBase" -> 0x0000000010000000L,
//+    "ResetVector" -> 0x80000000L,
//+    "MemMapBase" -> 0x0000000080000000L,
//     "MemMapRegionBits" -> 28,
//-    "MMIOBase" -> 0x00000000e0000000L,
//-    "MMIOSize" -> 0x0000000020000000L
//+    "MMIOBase" -> 0x0000000040600000L,
//+    "MMIOSize" -> 0x0000000001000000L
//   )
// }
// 
module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [8:0]  io_rreq_bits_setIdx,
  output [27:0] io_rresp_data_0_tag,
  output [1:0]  io_rresp_data_0__type,
  output [38:0] io_rresp_data_0_target,
  output [2:0]  io_rresp_data_0_brIdx,
  output        io_rresp_data_0_valid,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [27:0] io_wreq_bits_data_tag,
  input  [1:0]  io_wreq_bits_data__type,
  input  [38:0] io_wreq_bits_data_target,
  input  [2:0]  io_wreq_bits_data_brIdx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  reg  REG; // @[SRAMTemplate.scala 80:30]
  reg [8:0] value; // @[Counter.scala 60:40]
  wire  wrap_wrap = value == 9'h1ff; // @[Counter.scala 72:24]
  wire [8:0] _wrap_value_T_1 = value + 9'h1; // @[Counter.scala 76:24]
  wire  wrap = REG & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = wrap ? 1'h0 : REG; // @[SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  wire  _T = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
  wire [8:0] setIdx = REG ? value : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [72:0] _T_1 = {io_wreq_bits_data_tag,io_wreq_bits_data__type,io_wreq_bits_data_target,io_wreq_bits_data_brIdx
    ,1'h1}; // @[SRAMTemplate.scala 92:78]
  reg  REG_1; // @[Hold.scala 28:106]
  reg [72:0] r_0; // @[Reg.scala 27:20]
  wire [72:0] _GEN_14 = REG_1 ? array_RW0_rdata_0 : r_0; // @[Reg.scala 28:19 27:20 28:23]
  array array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_rdata_0(array_RW0_rdata_0)
  );
  assign io_rreq_ready = ~REG & _T; // @[SRAMTemplate.scala 101:33]
  assign io_rresp_data_0_tag = _GEN_14[72:45]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0__type = _GEN_14[44:43]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_target = _GEN_14[42:4]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_brIdx = _GEN_14[3:1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_valid = _GEN_14[0]; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = REG ? 73'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_en = realRen | wen;
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[Counter.scala 60:40]
      value <= 9'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      value <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    REG_1 <= io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
    if (reset) begin // @[Reg.scala 27:20]
      r_0 <= 73'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_0 <= array_RW0_rdata_0; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {3{`RANDOM}};
  r_0 = _RAND_3[72:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid,
  input  [38:0] io_in_pc_bits,
  output [38:0] io_out_target,
  output        io_out_valid,
  input         io_flush,
  output [2:0]  io_brIdx,
  output        io_crosslineJump,
  input         MOUFlushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[BPU.scala 302:19]
  wire  btb_reset; // @[BPU.scala 302:19]
  wire  btb_io_rreq_ready; // @[BPU.scala 302:19]
  wire  btb_io_rreq_valid; // @[BPU.scala 302:19]
  wire [8:0] btb_io_rreq_bits_setIdx; // @[BPU.scala 302:19]
  wire [27:0] btb_io_rresp_data_0_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_rresp_data_0__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_rresp_data_0_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_rresp_data_0_brIdx; // @[BPU.scala 302:19]
  wire  btb_io_rresp_data_0_valid; // @[BPU.scala 302:19]
  wire  btb_io_wreq_valid; // @[BPU.scala 302:19]
  wire [8:0] btb_io_wreq_bits_setIdx; // @[BPU.scala 302:19]
  wire [27:0] btb_io_wreq_bits_data_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_wreq_bits_data__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_wreq_bits_data_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_wreq_bits_data_brIdx; // @[BPU.scala 302:19]
  reg [1:0] pht [0:511]; // @[BPU.scala 336:16]
  wire  pht_MPORT_en; // @[BPU.scala 336:16]
  wire [8:0] pht_MPORT_addr; // @[BPU.scala 336:16]
  wire [1:0] pht_MPORT_data; // @[BPU.scala 336:16]
  wire  pht_MPORT_2_en; // @[BPU.scala 336:16]
  wire [8:0] pht_MPORT_2_addr; // @[BPU.scala 336:16]
  wire [1:0] pht_MPORT_2_data; // @[BPU.scala 336:16]
  wire [1:0] pht_MPORT_3_data; // @[BPU.scala 336:16]
  wire [8:0] pht_MPORT_3_addr; // @[BPU.scala 336:16]
  wire  pht_MPORT_3_mask; // @[BPU.scala 336:16]
  wire  pht_MPORT_3_en; // @[BPU.scala 336:16]
  reg [38:0] ras [0:15]; // @[BPU.scala 342:16]
  wire  ras_MPORT_1_en; // @[BPU.scala 342:16]
  wire [3:0] ras_MPORT_1_addr; // @[BPU.scala 342:16]
  wire [38:0] ras_MPORT_1_data; // @[BPU.scala 342:16]
  wire [38:0] ras_MPORT_4_data; // @[BPU.scala 342:16]
  wire [3:0] ras_MPORT_4_addr; // @[BPU.scala 342:16]
  wire  ras_MPORT_4_mask; // @[BPU.scala 342:16]
  wire  ras_MPORT_4_en; // @[BPU.scala 342:16]
  reg  flush; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = io_flush | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg [38:0] pcLatch; // @[Reg.scala 15:16]
  wire [27:0] btbRead_tag = btb_io_rresp_data_0_tag; // @[BPU.scala 315:21 316:11]
  wire  btbRead_valid = btb_io_rresp_data_0_valid; // @[BPU.scala 315:21 316:11]
  wire  _T_23 = btb_io_rreq_ready & btb_io_rreq_valid; // @[Decoupled.scala 40:37]
  reg  REG_1; // @[BPU.scala 320:93]
  wire [2:0] btbRead_brIdx = btb_io_rresp_data_0_brIdx; // @[BPU.scala 315:21 316:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:11] & ~flush & REG_1 & ~(pcLatch[1] & btbRead_brIdx[0]); // @[BPU.scala 320:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 327:40]
  reg  phtTaken; // @[Reg.scala 15:16]
  reg [3:0] value; // @[Counter.scala 60:40]
  reg [38:0] rasTarget; // @[Reg.scala 15:16]
  wire  _T_40 = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[BPU.scala 367:46]
  wire  _T_43 = ~bpuUpdateReq_pc[1]; // @[BPU.scala 367:72]
  wire [1:0] hi = {_T_40,bpuUpdateReq_pc[1]}; // @[Cat.scala 30:58]
  reg [1:0] cnt; // @[BPU.scala 389:20]
  reg  reqLatch_valid; // @[BPU.scala 390:25]
  reg [38:0] reqLatch_pc; // @[BPU.scala 390:25]
  reg  reqLatch_actualTaken; // @[BPU.scala 390:25]
  reg [6:0] reqLatch_fuOpType; // @[BPU.scala 390:25]
  wire  _T_53 = ~reqLatch_fuOpType[3]; // @[ALU.scala 63:30]
  wire  _T_54 = reqLatch_valid & _T_53; // @[BPU.scala 391:24]
  wire [1:0] _T_56 = cnt + 2'h1; // @[BPU.scala 393:33]
  wire [1:0] _T_58 = cnt - 2'h1; // @[BPU.scala 393:44]
  wire  _T_65 = reqLatch_actualTaken & cnt != 2'h3 | ~reqLatch_actualTaken & cnt != 2'h0; // @[BPU.scala 394:44]
  wire  _T_69 = bpuUpdateReq_fuOpType == 7'h5c; // @[BPU.scala 403:24]
  wire [3:0] _T_71 = value + 4'h1; // @[BPU.scala 404:26]
  wire [38:0] _T_73 = bpuUpdateReq_pc + 39'h2; // @[BPU.scala 404:55]
  wire [38:0] _T_75 = bpuUpdateReq_pc + 39'h4; // @[BPU.scala 404:69]
  wire  _T_78 = value == 4'h0; // @[BPU.scala 409:21]
  wire [3:0] _value_T_4 = value - 4'h1; // @[BPU.scala 412:53]
  wire [3:0] _value_T_5 = _T_78 ? 4'h0 : _value_T_4; // @[BPU.scala 412:22]
  wire [1:0] btbRead__type = btb_io_rresp_data_0__type; // @[BPU.scala 315:21 316:11]
  wire [38:0] btbRead_target = btb_io_rresp_data_0_target; // @[BPU.scala 315:21 316:11]
  wire [1:0] _T_82 = io_out_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_83 = {1'h1,crosslineJump,_T_82}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_28 = {{1'd0}, btbRead_brIdx}; // @[BPU.scala 419:30]
  wire [3:0] _T_84 = _GEN_28 & _T_83; // @[BPU.scala 419:30]
  wire  _T_88 = btbRead__type == 2'h0 ? phtTaken : rasTarget != 39'h0; // @[BPU.scala 420:32]
  SRAMTemplate btb ( // @[BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_rreq_ready(btb_io_rreq_ready),
    .io_rreq_valid(btb_io_rreq_valid),
    .io_rreq_bits_setIdx(btb_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(btb_io_rresp_data_0_tag),
    .io_rresp_data_0__type(btb_io_rresp_data_0__type),
    .io_rresp_data_0_target(btb_io_rresp_data_0_target),
    .io_rresp_data_0_brIdx(btb_io_rresp_data_0_brIdx),
    .io_rresp_data_0_valid(btb_io_rresp_data_0_valid),
    .io_wreq_valid(btb_io_wreq_valid),
    .io_wreq_bits_setIdx(btb_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(btb_io_wreq_bits_data_tag),
    .io_wreq_bits_data__type(btb_io_wreq_bits_data__type),
    .io_wreq_bits_data_target(btb_io_wreq_bits_data_target),
    .io_wreq_bits_data_brIdx(btb_io_wreq_bits_data_brIdx)
  );
  assign pht_MPORT_en = 1'h1;
  assign pht_MPORT_addr = io_in_pc_bits[10:2];
  assign pht_MPORT_data = pht[pht_MPORT_addr]; // @[BPU.scala 336:16]
  assign pht_MPORT_2_en = 1'h1;
  assign pht_MPORT_2_addr = bpuUpdateReq_pc[10:2];
  assign pht_MPORT_2_data = pht[pht_MPORT_2_addr]; // @[BPU.scala 336:16]
  assign pht_MPORT_3_data = reqLatch_actualTaken ? _T_56 : _T_58;
  assign pht_MPORT_3_addr = reqLatch_pc[10:2];
  assign pht_MPORT_3_mask = 1'h1;
  assign pht_MPORT_3_en = _T_54 & _T_65;
  assign ras_MPORT_1_en = 1'h1;
  assign ras_MPORT_1_addr = value;
  assign ras_MPORT_1_data = ras[ras_MPORT_1_addr]; // @[BPU.scala 342:16]
  assign ras_MPORT_4_data = bpuUpdateReq_isRVC ? _T_73 : _T_75;
  assign ras_MPORT_4_addr = value + 4'h1;
  assign ras_MPORT_4_mask = 1'h1;
  assign ras_MPORT_4_en = bpuUpdateReq_valid & _T_69;
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[BPU.scala 416:23]
  assign io_out_valid = btbHit & _T_88; // @[BPU.scala 420:26]
  assign io_brIdx = _T_84[2:0]; // @[BPU.scala 419:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 327:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[BPU.scala 308:29]
  assign btb_io_rreq_valid = io_in_pc_valid; // @[BPU.scala 311:22]
  assign btb_io_rreq_bits_setIdx = io_in_pc_bits[10:2]; // @[BPU.scala 35:65]
  assign btb_io_wreq_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[BPU.scala 375:43]
  assign btb_io_wreq_bits_setIdx = bpuUpdateReq_pc[10:2]; // @[BPU.scala 35:65]
  assign btb_io_wreq_bits_data_tag = bpuUpdateReq_pc[38:11]; // @[BPU.scala 35:65]
  assign btb_io_wreq_bits_data__type = bpuUpdateReq_btbType; // @[BPU.scala 377:26]
  assign btb_io_wreq_bits_data_target = bpuUpdateReq_actualTarget; // @[BPU.scala 377:26]
  assign btb_io_wreq_bits_data_brIdx = {hi,_T_43}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (pht_MPORT_3_en & pht_MPORT_3_mask) begin
      pht[pht_MPORT_3_addr] <= pht_MPORT_3_data; // @[BPU.scala 336:16]
    end
    if (ras_MPORT_4_en & ras_MPORT_4_mask) begin
      ras[ras_MPORT_4_addr] <= ras_MPORT_4_data; // @[BPU.scala 342:16]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      flush <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_1;
    end
    if (io_in_pc_valid) begin // @[Reg.scala 16:19]
      pcLatch <= io_in_pc_bits; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[BPU.scala 320:93]
      REG_1 <= 1'h0; // @[BPU.scala 320:93]
    end else begin
      REG_1 <= _T_23; // @[BPU.scala 320:93]
    end
    if (io_in_pc_valid) begin // @[Reg.scala 16:19]
      phtTaken <= pht_MPORT_data[1]; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 4'h0; // @[Counter.scala 60:40]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 403:45]
        value <= _T_71; // @[BPU.scala 406:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[BPU.scala 408:48]
        value <= _value_T_5; // @[BPU.scala 412:16]
      end
    end
    if (io_in_pc_valid) begin // @[Reg.scala 16:19]
      rasTarget <= ras_MPORT_1_data; // @[Reg.scala 16:23]
    end
    cnt <= pht_MPORT_2_data; // @[BPU.scala 389:20]
    reqLatch_valid <= bpuUpdateReq_valid; // @[BPU.scala 390:25]
    reqLatch_pc <= bpuUpdateReq_pc; // @[BPU.scala 390:25]
    reqLatch_actualTaken <= bpuUpdateReq_actualTaken; // @[BPU.scala 390:25]
    reqLatch_fuOpType <= bpuUpdateReq_fuOpType; // @[BPU.scala 390:25]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    pht[initvar] = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_1[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  flush = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  pcLatch = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  phtTaken = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[3:0];
  _RAND_7 = {2{`RANDOM}};
  rasTarget = _RAND_7[38:0];
  _RAND_8 = {1{`RANDOM}};
  cnt = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reqLatch_valid = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  reqLatch_pc = _RAND_10[38:0];
  _RAND_11 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_12[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [81:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [81:0] io_imem_resp_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input         flushICache,
  input         REG_0_valid,
  input  [38:0] REG_0_pc,
  input         REG_0_isMissPredict,
  input  [38:0] REG_0_actualTarget,
  input         REG_0_actualTaken,
  input  [6:0]  REG_0_fuOpType,
  input  [1:0]  REG_0_btbType,
  input         REG_0_isRVC,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[IFU.scala 326:19]
  wire  bp1_reset; // @[IFU.scala 326:19]
  wire  bp1_io_in_pc_valid; // @[IFU.scala 326:19]
  wire [38:0] bp1_io_in_pc_bits; // @[IFU.scala 326:19]
  wire [38:0] bp1_io_out_target; // @[IFU.scala 326:19]
  wire  bp1_io_out_valid; // @[IFU.scala 326:19]
  wire  bp1_io_flush; // @[IFU.scala 326:19]
  wire [2:0] bp1_io_brIdx; // @[IFU.scala 326:19]
  wire  bp1_io_crosslineJump; // @[IFU.scala 326:19]
  wire  bp1_MOUFlushICache; // @[IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_valid; // @[IFU.scala 326:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[IFU.scala 326:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[IFU.scala 326:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[IFU.scala 326:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[IFU.scala 326:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[IFU.scala 326:19]
  wire  bp1_MOUFlushTLB; // @[IFU.scala 326:19]
  reg [38:0] pc; // @[IFU.scala 322:19]
  wire  _T = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire  pcUpdate = io_redirect_valid | _T; // @[IFU.scala 323:36]
  wire [38:0] _T_3 = pc + 39'h2; // @[IFU.scala 324:28]
  wire [38:0] _T_5 = pc + 39'h4; // @[IFU.scala 324:38]
  wire [38:0] snpc = pc[1] ? _T_3 : _T_5; // @[IFU.scala 324:17]
  reg  crosslineJumpLatch; // @[IFU.scala 329:35]
  reg [38:0] crosslineJumpTarget; // @[Reg.scala 15:16]
  wire [38:0] pnpc = bp1_io_crosslineJump ? snpc : bp1_io_out_target; // @[IFU.scala 338:17]
  wire [38:0] _T_11 = bp1_io_out_valid ? pnpc : snpc; // @[IFU.scala 340:104]
  wire [38:0] _T_12 = crosslineJumpLatch ? crosslineJumpTarget : _T_11; // @[IFU.scala 340:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 340:16]
  wire  _T_13 = bp1_io_out_valid ? 1'h0 : 1'h1; // @[IFU.scala 341:114]
  wire  _T_15 = crosslineJumpLatch ? 1'h0 : bp1_io_crosslineJump | _T_13; // @[IFU.scala 341:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _T_15; // @[IFU.scala 341:21]
  wire [2:0] _T_16 = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[IFU.scala 349:29]
  wire [42:0] hi = {npcIsSeq,_T_16,npc}; // @[Cat.scala 30:58]
  wire  _T_34 = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | REG; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_35 = |io_flushVec; // @[IFU.scala 394:37]
  BPU_inorder bp1 ( // @[IFU.scala 326:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .MOUFlushICache(bp1_MOUFlushICache),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[IFU.scala 372:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[Cat.scala 30:58]
  assign io_imem_req_bits_user = {hi,pc}; // @[Cat.scala 30:58]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[IFU.scala 374:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[IFU.scala 391:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[IFU.scala 384:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[IFU.scala 386:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[IFU.scala 387:26]
  assign io_out_bits_exceptionVec_12 = io_ipf; // @[IFU.scala 390:44]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[IFU.scala 388:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[IFU.scala 367:21]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 340:16]
  assign bp1_io_flush = io_redirect_valid; // @[IFU.scala 358:16]
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_bpuUpdateReq_valid = REG_0_valid;
  assign bp1_bpuUpdateReq_pc = REG_0_pc;
  assign bp1_bpuUpdateReq_isMissPredict = REG_0_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = REG_0_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = REG_0_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = REG_0_fuOpType;
  assign bp1_bpuUpdateReq_btbType = REG_0_btbType;
  assign bp1_bpuUpdateReq_isRVC = REG_0_isRVC;
  assign bp1_MOUFlushTLB = flushTLB;
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 322:19]
      pc <= 39'h80000000; // @[IFU.scala 322:19]
    end else if (pcUpdate) begin // @[IFU.scala 360:19]
      if (io_redirect_valid) begin // @[IFU.scala 340:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[IFU.scala 340:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= _T_11;
      end
    end
    if (reset) begin // @[IFU.scala 329:35]
      crosslineJumpLatch <= 1'h0; // @[IFU.scala 329:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[IFU.scala 330:34]
      if (bp1_io_flush) begin // @[IFU.scala 331:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    if (bp1_io_crosslineJump) begin // @[Reg.scala 16:19]
      crosslineJumpTarget <= bp1_io_out_target; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_34) begin // @[StopWatch.scala 31:19]
      REG <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  REG = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  output        io_out_bits_crossPageIPFFix,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[NaiveIBF.scala 39:22]
  wire  _T_74 = state == 2'h2; // @[NaiveIBF.scala 90:23]
  wire  _T_75 = state == 2'h3; // @[NaiveIBF.scala 90:47]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[Cat.scala 30:58]
  reg [15:0] specialInstR; // @[NaiveIBF.scala 66:25]
  wire [31:0] _T_78 = {instIn[15:0],specialInstR}; // @[Cat.scala 30:58]
  wire  _T_1 = state == 2'h0; // @[NaiveIBF.scala 41:28]
  reg [2:0] pcOffsetR; // @[NaiveIBF.scala 40:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[NaiveIBF.scala 41:21]
  wire  _T_83 = 3'h0 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_87 = _T_83 ? instIn[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_84 = 3'h2 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_88 = _T_84 ? instIn[47:16] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_91 = _T_87 | _T_88; // @[Mux.scala 27:72]
  wire  _T_85 = 3'h4 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_89 = _T_85 ? instIn[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_92 = _T_91 | _T_89; // @[Mux.scala 27:72]
  wire  _T_86 = 3'h6 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_90 = _T_86 ? instIn[79:48] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_93 = _T_92 | _T_90; // @[Mux.scala 27:72]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _T_78 : _T_93; // @[NaiveIBF.scala 90:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[NaiveIBF.scala 34:26]
  wire  _T_3 = pcOffset == 3'h0; // @[NaiveIBF.scala 48:28]
  wire  _T_4 = ~isRVC; // @[NaiveIBF.scala 48:40]
  wire  _T_8 = pcOffset == 3'h4; // @[NaiveIBF.scala 48:72]
  wire  _T_14 = pcOffset == 3'h2; // @[NaiveIBF.scala 48:116]
  wire  _T_19 = pcOffset == 3'h6; // @[NaiveIBF.scala 48:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[NaiveIBF.scala 48:147]
  wire  _T_34 = _T_14 & _T_4; // @[NaiveIBF.scala 51:122]
  wire  _T_36 = ~io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:135]
  wire  rvcNext = _T_3 & (isRVC & ~io_in_bits_brIdx[0]) | _T_8 & (isRVC & ~io_in_bits_brIdx[0]) | _T_14 & _T_4 & ~
    io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:102]
  wire  _T_40 = _T_19 & _T_4; // @[NaiveIBF.scala 52:37]
  wire  rvcSpecial = _T_19 & _T_4 & ~io_in_bits_brIdx[2]; // @[NaiveIBF.scala 52:47]
  wire  rvcSpecialJump = _T_40 & io_in_bits_brIdx[2]; // @[NaiveIBF.scala 53:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[NaiveIBF.scala 54:24]
  wire  _T_49 = _T_1 | state == 2'h1; // @[NaiveIBF.scala 57:36]
  wire  flushIFU = (_T_1 | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[NaiveIBF.scala 57:87]
  wire  loadNextInstline = _T_49 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[NaiveIBF.scala 60:115]
  reg [38:0] specialPCR; // @[NaiveIBF.scala 64:23]
  reg [38:0] specialNPCR; // @[NaiveIBF.scala 65:24]
  reg  specialIPFR; // @[NaiveIBF.scala 67:28]
  wire  rvcForceLoadNext = _T_34 & io_in_bits_pnpc[2:0] == 3'h4 & _T_36; // @[NaiveIBF.scala 69:86]
  wire  _T_97 = rvcFinish | rvcNext; // @[NaiveIBF.scala 100:28]
  wire  _T_98 = rvcFinish | rvcForceLoadNext; // @[NaiveIBF.scala 101:28]
  wire [38:0] _T_100 = io_in_bits_pc + 39'h2; // @[NaiveIBF.scala 103:76]
  wire [38:0] _T_102 = io_in_bits_pc + 39'h4; // @[NaiveIBF.scala 103:95]
  wire [38:0] _T_103 = isRVC ? _T_100 : _T_102; // @[NaiveIBF.scala 103:55]
  wire [38:0] _T_104 = rvcFinish ? io_in_bits_pnpc : _T_103; // @[NaiveIBF.scala 103:23]
  wire  _T_105 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_0 = _T_105 & rvcFinish ? 2'h0 : state; // @[NaiveIBF.scala 104:{41,48} 39:22]
  wire [2:0] _T_109 = isRVC ? 3'h2 : 3'h4; // @[NaiveIBF.scala 107:38]
  wire [2:0] _T_111 = pcOffset + _T_109; // @[NaiveIBF.scala 107:33]
  wire [1:0] _GEN_1 = _T_105 & rvcNext ? 2'h1 : _GEN_0; // @[NaiveIBF.scala 105:39 106:17]
  wire [2:0] _GEN_2 = _T_105 & rvcNext ? _T_111 : pcOffsetR; // @[NaiveIBF.scala 105:39 107:21 40:26]
  wire [1:0] _GEN_3 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_1; // @[NaiveIBF.scala 109:40 110:17]
  wire [38:0] _T_121 = {io_in_bits_pc[38:3],pcOffsetR}; // @[Cat.scala 30:58]
  wire [38:0] _GEN_27 = 2'h3 == state ? specialPCR : 39'h0; // @[NaiveIBF.scala 161:15 98:18]
  wire [38:0] _GEN_32 = 2'h2 == state ? specialPCR : _GEN_27; // @[NaiveIBF.scala 149:15 98:18]
  wire [38:0] _GEN_40 = 2'h1 == state ? _T_121 : _GEN_32; // @[NaiveIBF.scala 126:15 98:18]
  wire [38:0] pcOut = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[NaiveIBF.scala 102:15 98:18]
  wire [38:0] _GEN_4 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[NaiveIBF.scala 109:40 111:22 64:23]
  wire [15:0] _GEN_5 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[NaiveIBF.scala 109:40 112:24 66:25]
  wire  _GEN_6 = rvcSpecial & io_in_valid ? io_in_bits_exceptionVec_12 : specialIPFR; // @[NaiveIBF.scala 109:40 113:23 67:28]
  wire [1:0] _GEN_7 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_3; // @[NaiveIBF.scala 115:44 116:17]
  wire [38:0] _GEN_8 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_4; // @[NaiveIBF.scala 115:44 117:22]
  wire [38:0] _GEN_9 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[NaiveIBF.scala 115:44 118:23 65:24]
  wire [15:0] _GEN_10 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_5; // @[NaiveIBF.scala 115:44 119:24]
  wire  _GEN_11 = rvcSpecialJump & io_in_valid ? io_in_bits_exceptionVec_12 : _GEN_6; // @[NaiveIBF.scala 115:44 120:23]
  wire [38:0] _T_123 = pcOut + 39'h2; // @[NaiveIBF.scala 127:68]
  wire [38:0] _T_125 = pcOut + 39'h4; // @[NaiveIBF.scala 127:79]
  wire [38:0] _T_126 = isRVC ? _T_123 : _T_125; // @[NaiveIBF.scala 127:55]
  wire [38:0] _T_127 = rvcFinish ? io_in_bits_pnpc : _T_126; // @[NaiveIBF.scala 127:23]
  wire [38:0] _T_141 = specialPCR + 39'h4; // @[NaiveIBF.scala 150:31]
  wire [1:0] _GEN_24 = _T_105 ? 2'h1 : state; // @[NaiveIBF.scala 154:28 155:17 39:22]
  wire [2:0] _GEN_25 = _T_105 ? 3'h2 : pcOffsetR; // @[NaiveIBF.scala 154:28 156:21 40:26]
  wire [1:0] _GEN_26 = _T_105 ? 2'h0 : state; // @[NaiveIBF.scala 166:28 167:17 39:22]
  wire [38:0] _GEN_28 = 2'h3 == state ? specialNPCR : 39'h0; // @[NaiveIBF.scala 162:17 98:18]
  wire  _GEN_29 = 2'h3 == state & io_in_valid; // @[NaiveIBF.scala 164:15 98:18]
  wire [1:0] _GEN_31 = 2'h3 == state ? _GEN_26 : state; // @[NaiveIBF.scala 98:18 39:22]
  wire [38:0] _GEN_33 = 2'h2 == state ? _T_141 : _GEN_28; // @[NaiveIBF.scala 150:17 98:18]
  wire  _GEN_34 = 2'h2 == state ? io_in_valid : _GEN_29; // @[NaiveIBF.scala 152:15 98:18]
  wire  _GEN_35 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[NaiveIBF.scala 153:15 98:18]
  wire [1:0] _GEN_36 = 2'h2 == state ? _GEN_24 : _GEN_31; // @[NaiveIBF.scala 98:18]
  wire [2:0] _GEN_37 = 2'h2 == state ? _GEN_25 : pcOffsetR; // @[NaiveIBF.scala 98:18 40:26]
  wire  _GEN_38 = 2'h1 == state ? _T_97 : _GEN_34; // @[NaiveIBF.scala 124:15 98:18]
  wire  _GEN_39 = 2'h1 == state ? _T_98 : _GEN_35; // @[NaiveIBF.scala 125:15 98:18]
  wire [38:0] _GEN_41 = 2'h1 == state ? _T_127 : _GEN_33; // @[NaiveIBF.scala 127:17 98:18]
  wire  canGo = 2'h0 == state ? rvcFinish | rvcNext : _GEN_38; // @[NaiveIBF.scala 100:15 98:18]
  wire  canIn = 2'h0 == state ? rvcFinish | rvcForceLoadNext : _GEN_39; // @[NaiveIBF.scala 101:15 98:18]
  wire [38:0] pnpcOut = 2'h0 == state ? _T_104 : _GEN_41; // @[NaiveIBF.scala 103:17 98:18]
  wire  _T_155 = pnpcOut == _T_125 & _T_4 | pnpcOut == _T_123 & isRVC ? 1'h0 : 1'h1; // @[NaiveIBF.scala 185:27]
  wire  _T_164 = _T_75 | _T_74; // @[NaiveIBF.scala 191:133]
  assign io_in_ready = ~io_in_valid | _T_105 & canIn | loadNextInstline; // @[NaiveIBF.scala 188:60]
  assign io_out_valid = io_in_valid & canGo; // @[NaiveIBF.scala 187:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[NaiveIBF.scala 184:21]
  assign io_out_bits_pc = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[NaiveIBF.scala 102:15 98:18]
  assign io_out_bits_pnpc = 2'h0 == state ? _T_104 : _GEN_41; // @[NaiveIBF.scala 103:17 98:18]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | specialIPFR & (_T_75 | _T_74); // @[NaiveIBF.scala 191:87]
  assign io_out_bits_brIdx = {{3'd0}, _T_155}; // @[NaiveIBF.scala 185:21]
  assign io_out_bits_crossPageIPFFix = io_in_bits_exceptionVec_12 & _T_164 & ~specialIPFR; // @[NaiveIBF.scala 192:130]
  always @(posedge clock) begin
    if (reset) begin // @[NaiveIBF.scala 39:22]
      state <= 2'h0; // @[NaiveIBF.scala 39:22]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else begin
        state <= _GEN_36;
      end
    end else begin
      state <= 2'h0; // @[NaiveIBF.scala 172:11]
    end
    if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 40:26]
      pcOffsetR <= 3'h0; // @[NaiveIBF.scala 40:26]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else begin
        pcOffsetR <= _GEN_37;
      end
    end
    if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end
    end
    if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 67:28]
      specialIPFR <= 1'h0; // @[NaiveIBF.scala 67:28]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[NaiveIBF.scala 98:18]
        specialIPFR <= _GEN_11;
      end else if (2'h1 == state) begin // @[NaiveIBF.scala 98:18]
        specialIPFR <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~flushIFU | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:59 assert(!flushIFU)\n"); // @[NaiveIBF.scala 59:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~flushIFU | reset)) begin
          $fatal; // @[NaiveIBF.scala 59:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  specialPCR = _RAND_3[38:0];
  _RAND_4 = {2{`RANDOM}};
  specialNPCR = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  specialIPFR = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decoder(
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_in_bits_crossPageIPFFix,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output        io_out_bits_ctrl_src1Type,
  output        io_out_bits_ctrl_src2Type,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output [4:0]  io_out_bits_ctrl_rfSrc1,
  output [4:0]  io_out_bits_ctrl_rfSrc2,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output [2:0]  io_out_bits_ctrl_vtag,
  output [4:0]  io_out_bits_ctrl_vec_addr,
  output [3:0]  io_out_bits_ctrl_length_k,
  output [1:0]  io_out_bits_ctrl_algorithm,
  output [63:0] io_out_bits_data_imm,
  output        io_isBranch,
  input         DTLBENABLE,
  input  [11:0] intrVecIDU
);
  wire [63:0] _T = io_in_bits_instr & 64'h707f; // @[Lookup.scala 31:38]
  wire  _T_1 = 64'h13 == _T; // @[Lookup.scala 31:38]
  wire [63:0] _T_2 = io_in_bits_instr & 64'hfc00707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 64'h1013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 64'h2013 == _T; // @[Lookup.scala 31:38]
  wire  _T_7 = 64'h3013 == _T; // @[Lookup.scala 31:38]
  wire  _T_9 = 64'h4013 == _T; // @[Lookup.scala 31:38]
  wire  _T_11 = 64'h5013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 64'h6013 == _T; // @[Lookup.scala 31:38]
  wire  _T_15 = 64'h7013 == _T; // @[Lookup.scala 31:38]
  wire  _T_17 = 64'h40005013 == _T_2; // @[Lookup.scala 31:38]
  wire [63:0] _T_18 = io_in_bits_instr & 64'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_19 = 64'h33 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_21 = 64'h1033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_23 = 64'h2033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_25 = 64'h3033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_27 = 64'h4033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_29 = 64'h5033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_31 = 64'h6033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_33 = 64'h7033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_35 = 64'h40000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_37 = 64'h40005033 == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_38 = io_in_bits_instr & 64'h7f; // @[Lookup.scala 31:38]
  wire  _T_39 = 64'h17 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_41 = 64'h37 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_43 = 64'h6f == _T_38; // @[Lookup.scala 31:38]
  wire  _T_45 = 64'h67 == _T; // @[Lookup.scala 31:38]
  wire  _T_47 = 64'h63 == _T; // @[Lookup.scala 31:38]
  wire  _T_49 = 64'h1063 == _T; // @[Lookup.scala 31:38]
  wire  _T_51 = 64'h4063 == _T; // @[Lookup.scala 31:38]
  wire  _T_53 = 64'h5063 == _T; // @[Lookup.scala 31:38]
  wire  _T_55 = 64'h6063 == _T; // @[Lookup.scala 31:38]
  wire  _T_57 = 64'h7063 == _T; // @[Lookup.scala 31:38]
  wire  _T_59 = 64'h3 == _T; // @[Lookup.scala 31:38]
  wire  _T_61 = 64'h1003 == _T; // @[Lookup.scala 31:38]
  wire  _T_63 = 64'h2003 == _T; // @[Lookup.scala 31:38]
  wire  _T_65 = 64'h4003 == _T; // @[Lookup.scala 31:38]
  wire  _T_67 = 64'h5003 == _T; // @[Lookup.scala 31:38]
  wire  _T_69 = 64'h23 == _T; // @[Lookup.scala 31:38]
  wire  _T_71 = 64'h1023 == _T; // @[Lookup.scala 31:38]
  wire  _T_73 = 64'h2023 == _T; // @[Lookup.scala 31:38]
  wire  _T_75 = 64'h1b == _T; // @[Lookup.scala 31:38]
  wire  _T_77 = 64'h101b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_79 = 64'h501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_81 = 64'h4000501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_83 = 64'h103b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_85 = 64'h503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_87 = 64'h4000503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_89 = 64'h3b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_91 = 64'h4000003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_93 = 64'h6003 == _T; // @[Lookup.scala 31:38]
  wire  _T_95 = 64'h3003 == _T; // @[Lookup.scala 31:38]
  wire  _T_97 = 64'h3023 == _T; // @[Lookup.scala 31:38]
  wire  _T_99 = 64'h6b == _T; // @[Lookup.scala 31:38]
  wire  _T_101 = 64'h2000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_103 = 64'h2001033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_105 = 64'h2002033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_107 = 64'h2003033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_109 = 64'h2004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_111 = 64'h2005033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_113 = 64'h2006033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_115 = 64'h2007033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_117 = 64'h200003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_119 = 64'h200403b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_121 = 64'h200503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_123 = 64'h200603b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_125 = 64'h200703b == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_126 = io_in_bits_instr & 64'hffffffff; // @[Lookup.scala 31:38]
  wire  _T_127 = 64'h0 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_128 = io_in_bits_instr & 64'he003; // @[Lookup.scala 31:38]
  wire  _T_129 = 64'h0 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_131 = 64'h4000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_133 = 64'h6000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_135 = 64'hc000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_137 = 64'he000 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_138 = io_in_bits_instr & 64'hef83; // @[Lookup.scala 31:38]
  wire  _T_139 = 64'h1 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_141 = 64'h1 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_143 = 64'h2001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_145 = 64'h4001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_147 = 64'h6101 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_149 = 64'h6001 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_150 = io_in_bits_instr & 64'hec03; // @[Lookup.scala 31:38]
  wire  _T_151 = 64'h8001 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_153 = 64'h8401 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_155 = 64'h8801 == _T_150; // @[Lookup.scala 31:38]
  wire [63:0] _T_156 = io_in_bits_instr & 64'hfc63; // @[Lookup.scala 31:38]
  wire  _T_157 = 64'h8c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_159 = 64'h8c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_161 = 64'h8c41 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_163 = 64'h8c61 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_165 = 64'h9c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_167 = 64'h9c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_169 = 64'ha001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_171 = 64'hc001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_173 = 64'he001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_175 = 64'h2 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_177 = 64'h4002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_179 = 64'h6002 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_180 = io_in_bits_instr & 64'hf07f; // @[Lookup.scala 31:38]
  wire  _T_181 = 64'h8002 == _T_180; // @[Lookup.scala 31:38]
  wire [63:0] _T_182 = io_in_bits_instr & 64'hf003; // @[Lookup.scala 31:38]
  wire  _T_183 = 64'h8002 == _T_182; // @[Lookup.scala 31:38]
  wire [63:0] _T_184 = io_in_bits_instr & 64'hffff; // @[Lookup.scala 31:38]
  wire  _T_185 = 64'h9002 == _T_184; // @[Lookup.scala 31:38]
  wire  _T_187 = 64'h9002 == _T_180; // @[Lookup.scala 31:38]
  wire  _T_189 = 64'h9002 == _T_182; // @[Lookup.scala 31:38]
  wire  _T_191 = 64'hc002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_193 = 64'he002 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_194 = io_in_bits_instr & 64'hff0ff07f; // @[Lookup.scala 31:38]
  wire  _T_195 = 64'h400b == _T_194; // @[Lookup.scala 31:38]
  wire [63:0] _T_196 = io_in_bits_instr & 64'hff0e707f; // @[Lookup.scala 31:38]
  wire  _T_197 = 64'h600b == _T_196; // @[Lookup.scala 31:38]
  wire  _T_199 = 64'h700b == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_200 = io_in_bits_instr & 64'hf800707f; // @[Lookup.scala 31:38]
  wire  _T_201 = 64'h200b == _T_200; // @[Lookup.scala 31:38]
  wire  _T_203 = 64'h300b == _T_200; // @[Lookup.scala 31:38]
  wire [63:0] _T_204 = io_in_bits_instr & 64'h7fff; // @[Lookup.scala 31:38]
  wire  _T_205 = 64'hb == _T_204; // @[Lookup.scala 31:38]
  wire  _T_207 = 64'h73 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_209 = 64'h100073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_211 = 64'h30200073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_213 = 64'hf == _T; // @[Lookup.scala 31:38]
  wire  _T_215 = 64'h10500073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_217 = 64'h10200073 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_218 = io_in_bits_instr & 64'hfe007fff; // @[Lookup.scala 31:38]
  wire  _T_219 = 64'h12000073 == _T_218; // @[Lookup.scala 31:38]
  wire [63:0] _T_220 = io_in_bits_instr & 64'hf9f0707f; // @[Lookup.scala 31:38]
  wire  _T_221 = 64'h1000302f == _T_220; // @[Lookup.scala 31:38]
  wire  _T_223 = 64'h1000202f == _T_220; // @[Lookup.scala 31:38]
  wire  _T_225 = 64'h1800302f == _T_200; // @[Lookup.scala 31:38]
  wire  _T_227 = 64'h1800202f == _T_200; // @[Lookup.scala 31:38]
  wire [63:0] _T_228 = io_in_bits_instr & 64'hf800607f; // @[Lookup.scala 31:38]
  wire  _T_229 = 64'h800202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_231 = 64'h202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_233 = 64'h2000202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_235 = 64'h6000202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_237 = 64'h4000202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_239 = 64'h8000202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_241 = 64'ha000202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_243 = 64'hc000202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_245 = 64'he000202f == _T_228; // @[Lookup.scala 31:38]
  wire  _T_247 = 64'h1073 == _T; // @[Lookup.scala 31:38]
  wire  _T_249 = 64'h2073 == _T; // @[Lookup.scala 31:38]
  wire  _T_251 = 64'h3073 == _T; // @[Lookup.scala 31:38]
  wire  _T_253 = 64'h5073 == _T; // @[Lookup.scala 31:38]
  wire  _T_255 = 64'h6073 == _T; // @[Lookup.scala 31:38]
  wire  _T_257 = 64'h7073 == _T; // @[Lookup.scala 31:38]
  wire  _T_259 = 64'h100f == _T_126; // @[Lookup.scala 31:38]
  wire [2:0] _T_261 = _T_257 ? 3'h4 : {{2'd0}, _T_259}; // @[Lookup.scala 33:37]
  wire [2:0] _T_262 = _T_255 ? 3'h4 : _T_261; // @[Lookup.scala 33:37]
  wire [2:0] _T_263 = _T_253 ? 3'h4 : _T_262; // @[Lookup.scala 33:37]
  wire [2:0] _T_264 = _T_251 ? 3'h4 : _T_263; // @[Lookup.scala 33:37]
  wire [2:0] _T_265 = _T_249 ? 3'h4 : _T_264; // @[Lookup.scala 33:37]
  wire [2:0] _T_266 = _T_247 ? 3'h4 : _T_265; // @[Lookup.scala 33:37]
  wire [2:0] _T_267 = _T_245 ? 3'h5 : _T_266; // @[Lookup.scala 33:37]
  wire [2:0] _T_268 = _T_243 ? 3'h5 : _T_267; // @[Lookup.scala 33:37]
  wire [2:0] _T_269 = _T_241 ? 3'h5 : _T_268; // @[Lookup.scala 33:37]
  wire [2:0] _T_270 = _T_239 ? 3'h5 : _T_269; // @[Lookup.scala 33:37]
  wire [2:0] _T_271 = _T_237 ? 3'h5 : _T_270; // @[Lookup.scala 33:37]
  wire [2:0] _T_272 = _T_235 ? 3'h5 : _T_271; // @[Lookup.scala 33:37]
  wire [2:0] _T_273 = _T_233 ? 3'h5 : _T_272; // @[Lookup.scala 33:37]
  wire [2:0] _T_274 = _T_231 ? 3'h5 : _T_273; // @[Lookup.scala 33:37]
  wire [2:0] _T_275 = _T_229 ? 3'h5 : _T_274; // @[Lookup.scala 33:37]
  wire [3:0] _T_276 = _T_227 ? 4'hf : {{1'd0}, _T_275}; // @[Lookup.scala 33:37]
  wire [3:0] _T_277 = _T_225 ? 4'hf : _T_276; // @[Lookup.scala 33:37]
  wire [3:0] _T_278 = _T_223 ? 4'h4 : _T_277; // @[Lookup.scala 33:37]
  wire [3:0] _T_279 = _T_221 ? 4'h4 : _T_278; // @[Lookup.scala 33:37]
  wire [3:0] _T_280 = _T_219 ? 4'h5 : _T_279; // @[Lookup.scala 33:37]
  wire [3:0] _T_281 = _T_217 ? 4'h4 : _T_280; // @[Lookup.scala 33:37]
  wire [3:0] _T_282 = _T_215 ? 4'h4 : _T_281; // @[Lookup.scala 33:37]
  wire [3:0] _T_283 = _T_213 ? 4'h2 : _T_282; // @[Lookup.scala 33:37]
  wire [3:0] _T_284 = _T_211 ? 4'h4 : _T_283; // @[Lookup.scala 33:37]
  wire [3:0] _T_285 = _T_209 ? 4'h4 : _T_284; // @[Lookup.scala 33:37]
  wire [3:0] _T_286 = _T_207 ? 4'h4 : _T_285; // @[Lookup.scala 33:37]
  wire [3:0] _T_287 = _T_205 ? 4'h4 : _T_286; // @[Lookup.scala 33:37]
  wire [3:0] _T_288 = _T_203 ? 4'h4 : _T_287; // @[Lookup.scala 33:37]
  wire [3:0] _T_289 = _T_201 ? 4'h4 : _T_288; // @[Lookup.scala 33:37]
  wire [3:0] _T_290 = _T_199 ? 4'h5 : _T_289; // @[Lookup.scala 33:37]
  wire [3:0] _T_291 = _T_197 ? 4'h6 : _T_290; // @[Lookup.scala 33:37]
  wire [3:0] _T_292 = _T_195 ? 4'h6 : _T_291; // @[Lookup.scala 33:37]
  wire [3:0] _T_293 = _T_193 ? 4'h2 : _T_292; // @[Lookup.scala 33:37]
  wire [3:0] _T_294 = _T_191 ? 4'h2 : _T_293; // @[Lookup.scala 33:37]
  wire [3:0] _T_295 = _T_189 ? 4'h5 : _T_294; // @[Lookup.scala 33:37]
  wire [3:0] _T_296 = _T_187 ? 4'h4 : _T_295; // @[Lookup.scala 33:37]
  wire [3:0] _T_297 = _T_185 ? 4'h4 : _T_296; // @[Lookup.scala 33:37]
  wire [3:0] _T_298 = _T_183 ? 4'h5 : _T_297; // @[Lookup.scala 33:37]
  wire [3:0] _T_299 = _T_181 ? 4'h4 : _T_298; // @[Lookup.scala 33:37]
  wire [3:0] _T_300 = _T_179 ? 4'h4 : _T_299; // @[Lookup.scala 33:37]
  wire [3:0] _T_301 = _T_177 ? 4'h4 : _T_300; // @[Lookup.scala 33:37]
  wire [3:0] _T_302 = _T_175 ? 4'h4 : _T_301; // @[Lookup.scala 33:37]
  wire [3:0] _T_303 = _T_173 ? 4'h1 : _T_302; // @[Lookup.scala 33:37]
  wire [3:0] _T_304 = _T_171 ? 4'h1 : _T_303; // @[Lookup.scala 33:37]
  wire [3:0] _T_305 = _T_169 ? 4'h7 : _T_304; // @[Lookup.scala 33:37]
  wire [3:0] _T_306 = _T_167 ? 4'h5 : _T_305; // @[Lookup.scala 33:37]
  wire [3:0] _T_307 = _T_165 ? 4'h5 : _T_306; // @[Lookup.scala 33:37]
  wire [3:0] _T_308 = _T_163 ? 4'h5 : _T_307; // @[Lookup.scala 33:37]
  wire [3:0] _T_309 = _T_161 ? 4'h5 : _T_308; // @[Lookup.scala 33:37]
  wire [3:0] _T_310 = _T_159 ? 4'h5 : _T_309; // @[Lookup.scala 33:37]
  wire [3:0] _T_311 = _T_157 ? 4'h5 : _T_310; // @[Lookup.scala 33:37]
  wire [3:0] _T_312 = _T_155 ? 4'h4 : _T_311; // @[Lookup.scala 33:37]
  wire [3:0] _T_313 = _T_153 ? 4'h4 : _T_312; // @[Lookup.scala 33:37]
  wire [3:0] _T_314 = _T_151 ? 4'h4 : _T_313; // @[Lookup.scala 33:37]
  wire [3:0] _T_315 = _T_149 ? 4'h4 : _T_314; // @[Lookup.scala 33:37]
  wire [3:0] _T_316 = _T_147 ? 4'h4 : _T_315; // @[Lookup.scala 33:37]
  wire [3:0] _T_317 = _T_145 ? 4'h4 : _T_316; // @[Lookup.scala 33:37]
  wire [3:0] _T_318 = _T_143 ? 4'h4 : _T_317; // @[Lookup.scala 33:37]
  wire [3:0] _T_319 = _T_141 ? 4'h4 : _T_318; // @[Lookup.scala 33:37]
  wire [3:0] _T_320 = _T_139 ? 4'h4 : _T_319; // @[Lookup.scala 33:37]
  wire [3:0] _T_321 = _T_137 ? 4'h2 : _T_320; // @[Lookup.scala 33:37]
  wire [3:0] _T_322 = _T_135 ? 4'h2 : _T_321; // @[Lookup.scala 33:37]
  wire [3:0] _T_323 = _T_133 ? 4'h4 : _T_322; // @[Lookup.scala 33:37]
  wire [3:0] _T_324 = _T_131 ? 4'h4 : _T_323; // @[Lookup.scala 33:37]
  wire [3:0] _T_325 = _T_129 ? 4'h4 : _T_324; // @[Lookup.scala 33:37]
  wire [3:0] _T_326 = _T_127 ? 4'h0 : _T_325; // @[Lookup.scala 33:37]
  wire [3:0] _T_327 = _T_125 ? 4'h5 : _T_326; // @[Lookup.scala 33:37]
  wire [3:0] _T_328 = _T_123 ? 4'h5 : _T_327; // @[Lookup.scala 33:37]
  wire [3:0] _T_329 = _T_121 ? 4'h5 : _T_328; // @[Lookup.scala 33:37]
  wire [3:0] _T_330 = _T_119 ? 4'h5 : _T_329; // @[Lookup.scala 33:37]
  wire [3:0] _T_331 = _T_117 ? 4'h5 : _T_330; // @[Lookup.scala 33:37]
  wire [3:0] _T_332 = _T_115 ? 4'h5 : _T_331; // @[Lookup.scala 33:37]
  wire [3:0] _T_333 = _T_113 ? 4'h5 : _T_332; // @[Lookup.scala 33:37]
  wire [3:0] _T_334 = _T_111 ? 4'h5 : _T_333; // @[Lookup.scala 33:37]
  wire [3:0] _T_335 = _T_109 ? 4'h5 : _T_334; // @[Lookup.scala 33:37]
  wire [3:0] _T_336 = _T_107 ? 4'h5 : _T_335; // @[Lookup.scala 33:37]
  wire [3:0] _T_337 = _T_105 ? 4'h5 : _T_336; // @[Lookup.scala 33:37]
  wire [3:0] _T_338 = _T_103 ? 4'h5 : _T_337; // @[Lookup.scala 33:37]
  wire [3:0] _T_339 = _T_101 ? 4'h5 : _T_338; // @[Lookup.scala 33:37]
  wire [3:0] _T_340 = _T_99 ? 4'h4 : _T_339; // @[Lookup.scala 33:37]
  wire [3:0] _T_341 = _T_97 ? 4'h2 : _T_340; // @[Lookup.scala 33:37]
  wire [3:0] _T_342 = _T_95 ? 4'h4 : _T_341; // @[Lookup.scala 33:37]
  wire [3:0] _T_343 = _T_93 ? 4'h4 : _T_342; // @[Lookup.scala 33:37]
  wire [3:0] _T_344 = _T_91 ? 4'h5 : _T_343; // @[Lookup.scala 33:37]
  wire [3:0] _T_345 = _T_89 ? 4'h5 : _T_344; // @[Lookup.scala 33:37]
  wire [3:0] _T_346 = _T_87 ? 4'h5 : _T_345; // @[Lookup.scala 33:37]
  wire [3:0] _T_347 = _T_85 ? 4'h5 : _T_346; // @[Lookup.scala 33:37]
  wire [3:0] _T_348 = _T_83 ? 4'h5 : _T_347; // @[Lookup.scala 33:37]
  wire [3:0] _T_349 = _T_81 ? 4'h4 : _T_348; // @[Lookup.scala 33:37]
  wire [3:0] _T_350 = _T_79 ? 4'h4 : _T_349; // @[Lookup.scala 33:37]
  wire [3:0] _T_351 = _T_77 ? 4'h4 : _T_350; // @[Lookup.scala 33:37]
  wire [3:0] _T_352 = _T_75 ? 4'h4 : _T_351; // @[Lookup.scala 33:37]
  wire [3:0] _T_353 = _T_73 ? 4'h2 : _T_352; // @[Lookup.scala 33:37]
  wire [3:0] _T_354 = _T_71 ? 4'h2 : _T_353; // @[Lookup.scala 33:37]
  wire [3:0] _T_355 = _T_69 ? 4'h2 : _T_354; // @[Lookup.scala 33:37]
  wire [3:0] _T_356 = _T_67 ? 4'h4 : _T_355; // @[Lookup.scala 33:37]
  wire [3:0] _T_357 = _T_65 ? 4'h4 : _T_356; // @[Lookup.scala 33:37]
  wire [3:0] _T_358 = _T_63 ? 4'h4 : _T_357; // @[Lookup.scala 33:37]
  wire [3:0] _T_359 = _T_61 ? 4'h4 : _T_358; // @[Lookup.scala 33:37]
  wire [3:0] _T_360 = _T_59 ? 4'h4 : _T_359; // @[Lookup.scala 33:37]
  wire [3:0] _T_361 = _T_57 ? 4'h1 : _T_360; // @[Lookup.scala 33:37]
  wire [3:0] _T_362 = _T_55 ? 4'h1 : _T_361; // @[Lookup.scala 33:37]
  wire [3:0] _T_363 = _T_53 ? 4'h1 : _T_362; // @[Lookup.scala 33:37]
  wire [3:0] _T_364 = _T_51 ? 4'h1 : _T_363; // @[Lookup.scala 33:37]
  wire [3:0] _T_365 = _T_49 ? 4'h1 : _T_364; // @[Lookup.scala 33:37]
  wire [3:0] _T_366 = _T_47 ? 4'h1 : _T_365; // @[Lookup.scala 33:37]
  wire [3:0] _T_367 = _T_45 ? 4'h4 : _T_366; // @[Lookup.scala 33:37]
  wire [3:0] _T_368 = _T_43 ? 4'h7 : _T_367; // @[Lookup.scala 33:37]
  wire [3:0] _T_369 = _T_41 ? 4'h6 : _T_368; // @[Lookup.scala 33:37]
  wire [3:0] _T_370 = _T_39 ? 4'h6 : _T_369; // @[Lookup.scala 33:37]
  wire [3:0] _T_371 = _T_37 ? 4'h5 : _T_370; // @[Lookup.scala 33:37]
  wire [3:0] _T_372 = _T_35 ? 4'h5 : _T_371; // @[Lookup.scala 33:37]
  wire [3:0] _T_373 = _T_33 ? 4'h5 : _T_372; // @[Lookup.scala 33:37]
  wire [3:0] _T_374 = _T_31 ? 4'h5 : _T_373; // @[Lookup.scala 33:37]
  wire [3:0] _T_375 = _T_29 ? 4'h5 : _T_374; // @[Lookup.scala 33:37]
  wire [3:0] _T_376 = _T_27 ? 4'h5 : _T_375; // @[Lookup.scala 33:37]
  wire [3:0] _T_377 = _T_25 ? 4'h5 : _T_376; // @[Lookup.scala 33:37]
  wire [3:0] _T_378 = _T_23 ? 4'h5 : _T_377; // @[Lookup.scala 33:37]
  wire [3:0] _T_379 = _T_21 ? 4'h5 : _T_378; // @[Lookup.scala 33:37]
  wire [3:0] _T_380 = _T_19 ? 4'h5 : _T_379; // @[Lookup.scala 33:37]
  wire [3:0] _T_381 = _T_17 ? 4'h4 : _T_380; // @[Lookup.scala 33:37]
  wire [3:0] _T_382 = _T_15 ? 4'h4 : _T_381; // @[Lookup.scala 33:37]
  wire [3:0] _T_383 = _T_13 ? 4'h4 : _T_382; // @[Lookup.scala 33:37]
  wire [3:0] _T_384 = _T_11 ? 4'h4 : _T_383; // @[Lookup.scala 33:37]
  wire [3:0] _T_385 = _T_9 ? 4'h4 : _T_384; // @[Lookup.scala 33:37]
  wire [3:0] _T_386 = _T_7 ? 4'h4 : _T_385; // @[Lookup.scala 33:37]
  wire [3:0] _T_387 = _T_5 ? 4'h4 : _T_386; // @[Lookup.scala 33:37]
  wire [3:0] _T_388 = _T_3 ? 4'h4 : _T_387; // @[Lookup.scala 33:37]
  wire [3:0] decodeList_0 = _T_1 ? 4'h4 : _T_388; // @[Lookup.scala 33:37]
  wire [2:0] _T_389 = _T_259 ? 3'h4 : 3'h3; // @[Lookup.scala 33:37]
  wire [2:0] _T_390 = _T_257 ? 3'h3 : _T_389; // @[Lookup.scala 33:37]
  wire [2:0] _T_391 = _T_255 ? 3'h3 : _T_390; // @[Lookup.scala 33:37]
  wire [2:0] _T_392 = _T_253 ? 3'h3 : _T_391; // @[Lookup.scala 33:37]
  wire [2:0] _T_393 = _T_251 ? 3'h3 : _T_392; // @[Lookup.scala 33:37]
  wire [2:0] _T_394 = _T_249 ? 3'h3 : _T_393; // @[Lookup.scala 33:37]
  wire [2:0] _T_395 = _T_247 ? 3'h3 : _T_394; // @[Lookup.scala 33:37]
  wire [2:0] _T_396 = _T_245 ? 3'h1 : _T_395; // @[Lookup.scala 33:37]
  wire [2:0] _T_397 = _T_243 ? 3'h1 : _T_396; // @[Lookup.scala 33:37]
  wire [2:0] _T_398 = _T_241 ? 3'h1 : _T_397; // @[Lookup.scala 33:37]
  wire [2:0] _T_399 = _T_239 ? 3'h1 : _T_398; // @[Lookup.scala 33:37]
  wire [2:0] _T_400 = _T_237 ? 3'h1 : _T_399; // @[Lookup.scala 33:37]
  wire [2:0] _T_401 = _T_235 ? 3'h1 : _T_400; // @[Lookup.scala 33:37]
  wire [2:0] _T_402 = _T_233 ? 3'h1 : _T_401; // @[Lookup.scala 33:37]
  wire [2:0] _T_403 = _T_231 ? 3'h1 : _T_402; // @[Lookup.scala 33:37]
  wire [2:0] _T_404 = _T_229 ? 3'h1 : _T_403; // @[Lookup.scala 33:37]
  wire [2:0] _T_405 = _T_227 ? 3'h1 : _T_404; // @[Lookup.scala 33:37]
  wire [2:0] _T_406 = _T_225 ? 3'h1 : _T_405; // @[Lookup.scala 33:37]
  wire [2:0] _T_407 = _T_223 ? 3'h1 : _T_406; // @[Lookup.scala 33:37]
  wire [2:0] _T_408 = _T_221 ? 3'h1 : _T_407; // @[Lookup.scala 33:37]
  wire [2:0] _T_409 = _T_219 ? 3'h4 : _T_408; // @[Lookup.scala 33:37]
  wire [2:0] _T_410 = _T_217 ? 3'h3 : _T_409; // @[Lookup.scala 33:37]
  wire [2:0] _T_411 = _T_215 ? 3'h0 : _T_410; // @[Lookup.scala 33:37]
  wire [2:0] _T_412 = _T_213 ? 3'h4 : _T_411; // @[Lookup.scala 33:37]
  wire [2:0] _T_413 = _T_211 ? 3'h3 : _T_412; // @[Lookup.scala 33:37]
  wire [2:0] _T_414 = _T_209 ? 3'h3 : _T_413; // @[Lookup.scala 33:37]
  wire [2:0] _T_415 = _T_207 ? 3'h3 : _T_414; // @[Lookup.scala 33:37]
  wire [2:0] _T_416 = _T_205 ? 3'h5 : _T_415; // @[Lookup.scala 33:37]
  wire [2:0] _T_417 = _T_203 ? 3'h5 : _T_416; // @[Lookup.scala 33:37]
  wire [2:0] _T_418 = _T_201 ? 3'h5 : _T_417; // @[Lookup.scala 33:37]
  wire [2:0] _T_419 = _T_199 ? 3'h5 : _T_418; // @[Lookup.scala 33:37]
  wire [2:0] _T_420 = _T_197 ? 3'h5 : _T_419; // @[Lookup.scala 33:37]
  wire [2:0] _T_421 = _T_195 ? 3'h5 : _T_420; // @[Lookup.scala 33:37]
  wire [2:0] _T_422 = _T_193 ? 3'h1 : _T_421; // @[Lookup.scala 33:37]
  wire [2:0] _T_423 = _T_191 ? 3'h1 : _T_422; // @[Lookup.scala 33:37]
  wire [2:0] _T_424 = _T_189 ? 3'h0 : _T_423; // @[Lookup.scala 33:37]
  wire [2:0] _T_425 = _T_187 ? 3'h0 : _T_424; // @[Lookup.scala 33:37]
  wire [2:0] _T_426 = _T_185 ? 3'h3 : _T_425; // @[Lookup.scala 33:37]
  wire [2:0] _T_427 = _T_183 ? 3'h0 : _T_426; // @[Lookup.scala 33:37]
  wire [2:0] _T_428 = _T_181 ? 3'h0 : _T_427; // @[Lookup.scala 33:37]
  wire [2:0] _T_429 = _T_179 ? 3'h1 : _T_428; // @[Lookup.scala 33:37]
  wire [2:0] _T_430 = _T_177 ? 3'h1 : _T_429; // @[Lookup.scala 33:37]
  wire [2:0] _T_431 = _T_175 ? 3'h0 : _T_430; // @[Lookup.scala 33:37]
  wire [2:0] _T_432 = _T_173 ? 3'h0 : _T_431; // @[Lookup.scala 33:37]
  wire [2:0] _T_433 = _T_171 ? 3'h0 : _T_432; // @[Lookup.scala 33:37]
  wire [2:0] _T_434 = _T_169 ? 3'h0 : _T_433; // @[Lookup.scala 33:37]
  wire [2:0] _T_435 = _T_167 ? 3'h0 : _T_434; // @[Lookup.scala 33:37]
  wire [2:0] _T_436 = _T_165 ? 3'h0 : _T_435; // @[Lookup.scala 33:37]
  wire [2:0] _T_437 = _T_163 ? 3'h0 : _T_436; // @[Lookup.scala 33:37]
  wire [2:0] _T_438 = _T_161 ? 3'h0 : _T_437; // @[Lookup.scala 33:37]
  wire [2:0] _T_439 = _T_159 ? 3'h0 : _T_438; // @[Lookup.scala 33:37]
  wire [2:0] _T_440 = _T_157 ? 3'h0 : _T_439; // @[Lookup.scala 33:37]
  wire [2:0] _T_441 = _T_155 ? 3'h0 : _T_440; // @[Lookup.scala 33:37]
  wire [2:0] _T_442 = _T_153 ? 3'h0 : _T_441; // @[Lookup.scala 33:37]
  wire [2:0] _T_443 = _T_151 ? 3'h0 : _T_442; // @[Lookup.scala 33:37]
  wire [2:0] _T_444 = _T_149 ? 3'h0 : _T_443; // @[Lookup.scala 33:37]
  wire [2:0] _T_445 = _T_147 ? 3'h0 : _T_444; // @[Lookup.scala 33:37]
  wire [2:0] _T_446 = _T_145 ? 3'h0 : _T_445; // @[Lookup.scala 33:37]
  wire [2:0] _T_447 = _T_143 ? 3'h0 : _T_446; // @[Lookup.scala 33:37]
  wire [2:0] _T_448 = _T_141 ? 3'h0 : _T_447; // @[Lookup.scala 33:37]
  wire [2:0] _T_449 = _T_139 ? 3'h0 : _T_448; // @[Lookup.scala 33:37]
  wire [2:0] _T_450 = _T_137 ? 3'h1 : _T_449; // @[Lookup.scala 33:37]
  wire [2:0] _T_451 = _T_135 ? 3'h1 : _T_450; // @[Lookup.scala 33:37]
  wire [2:0] _T_452 = _T_133 ? 3'h1 : _T_451; // @[Lookup.scala 33:37]
  wire [2:0] _T_453 = _T_131 ? 3'h1 : _T_452; // @[Lookup.scala 33:37]
  wire [2:0] _T_454 = _T_129 ? 3'h0 : _T_453; // @[Lookup.scala 33:37]
  wire [2:0] _T_455 = _T_127 ? 3'h3 : _T_454; // @[Lookup.scala 33:37]
  wire [2:0] _T_456 = _T_125 ? 3'h2 : _T_455; // @[Lookup.scala 33:37]
  wire [2:0] _T_457 = _T_123 ? 3'h2 : _T_456; // @[Lookup.scala 33:37]
  wire [2:0] _T_458 = _T_121 ? 3'h2 : _T_457; // @[Lookup.scala 33:37]
  wire [2:0] _T_459 = _T_119 ? 3'h2 : _T_458; // @[Lookup.scala 33:37]
  wire [2:0] _T_460 = _T_117 ? 3'h2 : _T_459; // @[Lookup.scala 33:37]
  wire [2:0] _T_461 = _T_115 ? 3'h2 : _T_460; // @[Lookup.scala 33:37]
  wire [2:0] _T_462 = _T_113 ? 3'h2 : _T_461; // @[Lookup.scala 33:37]
  wire [2:0] _T_463 = _T_111 ? 3'h2 : _T_462; // @[Lookup.scala 33:37]
  wire [2:0] _T_464 = _T_109 ? 3'h2 : _T_463; // @[Lookup.scala 33:37]
  wire [2:0] _T_465 = _T_107 ? 3'h2 : _T_464; // @[Lookup.scala 33:37]
  wire [2:0] _T_466 = _T_105 ? 3'h2 : _T_465; // @[Lookup.scala 33:37]
  wire [2:0] _T_467 = _T_103 ? 3'h2 : _T_466; // @[Lookup.scala 33:37]
  wire [2:0] _T_468 = _T_101 ? 3'h2 : _T_467; // @[Lookup.scala 33:37]
  wire [2:0] _T_469 = _T_99 ? 3'h3 : _T_468; // @[Lookup.scala 33:37]
  wire [2:0] _T_470 = _T_97 ? 3'h1 : _T_469; // @[Lookup.scala 33:37]
  wire [2:0] _T_471 = _T_95 ? 3'h1 : _T_470; // @[Lookup.scala 33:37]
  wire [2:0] _T_472 = _T_93 ? 3'h1 : _T_471; // @[Lookup.scala 33:37]
  wire [2:0] _T_473 = _T_91 ? 3'h0 : _T_472; // @[Lookup.scala 33:37]
  wire [2:0] _T_474 = _T_89 ? 3'h0 : _T_473; // @[Lookup.scala 33:37]
  wire [2:0] _T_475 = _T_87 ? 3'h0 : _T_474; // @[Lookup.scala 33:37]
  wire [2:0] _T_476 = _T_85 ? 3'h0 : _T_475; // @[Lookup.scala 33:37]
  wire [2:0] _T_477 = _T_83 ? 3'h0 : _T_476; // @[Lookup.scala 33:37]
  wire [2:0] _T_478 = _T_81 ? 3'h0 : _T_477; // @[Lookup.scala 33:37]
  wire [2:0] _T_479 = _T_79 ? 3'h0 : _T_478; // @[Lookup.scala 33:37]
  wire [2:0] _T_480 = _T_77 ? 3'h0 : _T_479; // @[Lookup.scala 33:37]
  wire [2:0] _T_481 = _T_75 ? 3'h0 : _T_480; // @[Lookup.scala 33:37]
  wire [2:0] _T_482 = _T_73 ? 3'h1 : _T_481; // @[Lookup.scala 33:37]
  wire [2:0] _T_483 = _T_71 ? 3'h1 : _T_482; // @[Lookup.scala 33:37]
  wire [2:0] _T_484 = _T_69 ? 3'h1 : _T_483; // @[Lookup.scala 33:37]
  wire [2:0] _T_485 = _T_67 ? 3'h1 : _T_484; // @[Lookup.scala 33:37]
  wire [2:0] _T_486 = _T_65 ? 3'h1 : _T_485; // @[Lookup.scala 33:37]
  wire [2:0] _T_487 = _T_63 ? 3'h1 : _T_486; // @[Lookup.scala 33:37]
  wire [2:0] _T_488 = _T_61 ? 3'h1 : _T_487; // @[Lookup.scala 33:37]
  wire [2:0] _T_489 = _T_59 ? 3'h1 : _T_488; // @[Lookup.scala 33:37]
  wire [2:0] _T_490 = _T_57 ? 3'h0 : _T_489; // @[Lookup.scala 33:37]
  wire [2:0] _T_491 = _T_55 ? 3'h0 : _T_490; // @[Lookup.scala 33:37]
  wire [2:0] _T_492 = _T_53 ? 3'h0 : _T_491; // @[Lookup.scala 33:37]
  wire [2:0] _T_493 = _T_51 ? 3'h0 : _T_492; // @[Lookup.scala 33:37]
  wire [2:0] _T_494 = _T_49 ? 3'h0 : _T_493; // @[Lookup.scala 33:37]
  wire [2:0] _T_495 = _T_47 ? 3'h0 : _T_494; // @[Lookup.scala 33:37]
  wire [2:0] _T_496 = _T_45 ? 3'h0 : _T_495; // @[Lookup.scala 33:37]
  wire [2:0] _T_497 = _T_43 ? 3'h0 : _T_496; // @[Lookup.scala 33:37]
  wire [2:0] _T_498 = _T_41 ? 3'h0 : _T_497; // @[Lookup.scala 33:37]
  wire [2:0] _T_499 = _T_39 ? 3'h0 : _T_498; // @[Lookup.scala 33:37]
  wire [2:0] _T_500 = _T_37 ? 3'h0 : _T_499; // @[Lookup.scala 33:37]
  wire [2:0] _T_501 = _T_35 ? 3'h0 : _T_500; // @[Lookup.scala 33:37]
  wire [2:0] _T_502 = _T_33 ? 3'h0 : _T_501; // @[Lookup.scala 33:37]
  wire [2:0] _T_503 = _T_31 ? 3'h0 : _T_502; // @[Lookup.scala 33:37]
  wire [2:0] _T_504 = _T_29 ? 3'h0 : _T_503; // @[Lookup.scala 33:37]
  wire [2:0] _T_505 = _T_27 ? 3'h0 : _T_504; // @[Lookup.scala 33:37]
  wire [2:0] _T_506 = _T_25 ? 3'h0 : _T_505; // @[Lookup.scala 33:37]
  wire [2:0] _T_507 = _T_23 ? 3'h0 : _T_506; // @[Lookup.scala 33:37]
  wire [2:0] _T_508 = _T_21 ? 3'h0 : _T_507; // @[Lookup.scala 33:37]
  wire [2:0] _T_509 = _T_19 ? 3'h0 : _T_508; // @[Lookup.scala 33:37]
  wire [2:0] _T_510 = _T_17 ? 3'h0 : _T_509; // @[Lookup.scala 33:37]
  wire [2:0] _T_511 = _T_15 ? 3'h0 : _T_510; // @[Lookup.scala 33:37]
  wire [2:0] _T_512 = _T_13 ? 3'h0 : _T_511; // @[Lookup.scala 33:37]
  wire [2:0] _T_513 = _T_11 ? 3'h0 : _T_512; // @[Lookup.scala 33:37]
  wire [2:0] _T_514 = _T_9 ? 3'h0 : _T_513; // @[Lookup.scala 33:37]
  wire [2:0] _T_515 = _T_7 ? 3'h0 : _T_514; // @[Lookup.scala 33:37]
  wire [2:0] _T_516 = _T_5 ? 3'h0 : _T_515; // @[Lookup.scala 33:37]
  wire [2:0] _T_517 = _T_3 ? 3'h0 : _T_516; // @[Lookup.scala 33:37]
  wire [2:0] decodeList_1 = _T_1 ? 3'h0 : _T_517; // @[Lookup.scala 33:37]
  wire [2:0] _T_519 = _T_257 ? 3'h7 : {{2'd0}, _T_259}; // @[Lookup.scala 33:37]
  wire [2:0] _T_520 = _T_255 ? 3'h6 : _T_519; // @[Lookup.scala 33:37]
  wire [2:0] _T_521 = _T_253 ? 3'h5 : _T_520; // @[Lookup.scala 33:37]
  wire [2:0] _T_522 = _T_251 ? 3'h3 : _T_521; // @[Lookup.scala 33:37]
  wire [2:0] _T_523 = _T_249 ? 3'h2 : _T_522; // @[Lookup.scala 33:37]
  wire [2:0] _T_524 = _T_247 ? 3'h1 : _T_523; // @[Lookup.scala 33:37]
  wire [5:0] _T_525 = _T_245 ? 6'h32 : {{3'd0}, _T_524}; // @[Lookup.scala 33:37]
  wire [5:0] _T_526 = _T_243 ? 6'h31 : _T_525; // @[Lookup.scala 33:37]
  wire [5:0] _T_527 = _T_241 ? 6'h30 : _T_526; // @[Lookup.scala 33:37]
  wire [5:0] _T_528 = _T_239 ? 6'h37 : _T_527; // @[Lookup.scala 33:37]
  wire [5:0] _T_529 = _T_237 ? 6'h26 : _T_528; // @[Lookup.scala 33:37]
  wire [5:0] _T_530 = _T_235 ? 6'h25 : _T_529; // @[Lookup.scala 33:37]
  wire [5:0] _T_531 = _T_233 ? 6'h24 : _T_530; // @[Lookup.scala 33:37]
  wire [6:0] _T_532 = _T_231 ? 7'h63 : {{1'd0}, _T_531}; // @[Lookup.scala 33:37]
  wire [6:0] _T_533 = _T_229 ? 7'h22 : _T_532; // @[Lookup.scala 33:37]
  wire [6:0] _T_534 = _T_227 ? 7'h21 : _T_533; // @[Lookup.scala 33:37]
  wire [6:0] _T_535 = _T_225 ? 7'h21 : _T_534; // @[Lookup.scala 33:37]
  wire [6:0] _T_536 = _T_223 ? 7'h20 : _T_535; // @[Lookup.scala 33:37]
  wire [6:0] _T_537 = _T_221 ? 7'h20 : _T_536; // @[Lookup.scala 33:37]
  wire [6:0] _T_538 = _T_219 ? 7'h2 : _T_537; // @[Lookup.scala 33:37]
  wire [6:0] _T_539 = _T_217 ? 7'h0 : _T_538; // @[Lookup.scala 33:37]
  wire [6:0] _T_540 = _T_215 ? 7'h40 : _T_539; // @[Lookup.scala 33:37]
  wire [6:0] _T_541 = _T_213 ? 7'h0 : _T_540; // @[Lookup.scala 33:37]
  wire [6:0] _T_542 = _T_211 ? 7'h0 : _T_541; // @[Lookup.scala 33:37]
  wire [6:0] _T_543 = _T_209 ? 7'h0 : _T_542; // @[Lookup.scala 33:37]
  wire [6:0] _T_544 = _T_207 ? 7'h0 : _T_543; // @[Lookup.scala 33:37]
  wire [6:0] _T_545 = _T_205 ? 7'h9 : _T_544; // @[Lookup.scala 33:37]
  wire [6:0] _T_546 = _T_203 ? 7'ha : _T_545; // @[Lookup.scala 33:37]
  wire [6:0] _T_547 = _T_201 ? 7'hc : _T_546; // @[Lookup.scala 33:37]
  wire [6:0] _T_548 = _T_199 ? 7'h4 : _T_547; // @[Lookup.scala 33:37]
  wire [6:0] _T_549 = _T_197 ? 7'h2 : _T_548; // @[Lookup.scala 33:37]
  wire [6:0] _T_550 = _T_195 ? 7'h1 : _T_549; // @[Lookup.scala 33:37]
  wire [6:0] _T_551 = _T_193 ? 7'hb : _T_550; // @[Lookup.scala 33:37]
  wire [6:0] _T_552 = _T_191 ? 7'ha : _T_551; // @[Lookup.scala 33:37]
  wire [6:0] _T_553 = _T_189 ? 7'h40 : _T_552; // @[Lookup.scala 33:37]
  wire [6:0] _T_554 = _T_187 ? 7'h5a : _T_553; // @[Lookup.scala 33:37]
  wire [6:0] _T_555 = _T_185 ? 7'h0 : _T_554; // @[Lookup.scala 33:37]
  wire [6:0] _T_556 = _T_183 ? 7'h40 : _T_555; // @[Lookup.scala 33:37]
  wire [6:0] _T_557 = _T_181 ? 7'h5a : _T_556; // @[Lookup.scala 33:37]
  wire [6:0] _T_558 = _T_179 ? 7'h3 : _T_557; // @[Lookup.scala 33:37]
  wire [6:0] _T_559 = _T_177 ? 7'h2 : _T_558; // @[Lookup.scala 33:37]
  wire [6:0] _T_560 = _T_175 ? 7'h1 : _T_559; // @[Lookup.scala 33:37]
  wire [6:0] _T_561 = _T_173 ? 7'h11 : _T_560; // @[Lookup.scala 33:37]
  wire [6:0] _T_562 = _T_171 ? 7'h10 : _T_561; // @[Lookup.scala 33:37]
  wire [6:0] _T_563 = _T_169 ? 7'h58 : _T_562; // @[Lookup.scala 33:37]
  wire [6:0] _T_564 = _T_167 ? 7'h60 : _T_563; // @[Lookup.scala 33:37]
  wire [6:0] _T_565 = _T_165 ? 7'h28 : _T_564; // @[Lookup.scala 33:37]
  wire [6:0] _T_566 = _T_163 ? 7'h7 : _T_565; // @[Lookup.scala 33:37]
  wire [6:0] _T_567 = _T_161 ? 7'h6 : _T_566; // @[Lookup.scala 33:37]
  wire [6:0] _T_568 = _T_159 ? 7'h4 : _T_567; // @[Lookup.scala 33:37]
  wire [6:0] _T_569 = _T_157 ? 7'h8 : _T_568; // @[Lookup.scala 33:37]
  wire [6:0] _T_570 = _T_155 ? 7'h7 : _T_569; // @[Lookup.scala 33:37]
  wire [6:0] _T_571 = _T_153 ? 7'hd : _T_570; // @[Lookup.scala 33:37]
  wire [6:0] _T_572 = _T_151 ? 7'h5 : _T_571; // @[Lookup.scala 33:37]
  wire [6:0] _T_573 = _T_149 ? 7'h40 : _T_572; // @[Lookup.scala 33:37]
  wire [6:0] _T_574 = _T_147 ? 7'h40 : _T_573; // @[Lookup.scala 33:37]
  wire [6:0] _T_575 = _T_145 ? 7'h40 : _T_574; // @[Lookup.scala 33:37]
  wire [6:0] _T_576 = _T_143 ? 7'h60 : _T_575; // @[Lookup.scala 33:37]
  wire [6:0] _T_577 = _T_141 ? 7'h40 : _T_576; // @[Lookup.scala 33:37]
  wire [6:0] _T_578 = _T_139 ? 7'h40 : _T_577; // @[Lookup.scala 33:37]
  wire [6:0] _T_579 = _T_137 ? 7'hb : _T_578; // @[Lookup.scala 33:37]
  wire [6:0] _T_580 = _T_135 ? 7'ha : _T_579; // @[Lookup.scala 33:37]
  wire [6:0] _T_581 = _T_133 ? 7'h3 : _T_580; // @[Lookup.scala 33:37]
  wire [6:0] _T_582 = _T_131 ? 7'h2 : _T_581; // @[Lookup.scala 33:37]
  wire [6:0] _T_583 = _T_129 ? 7'h40 : _T_582; // @[Lookup.scala 33:37]
  wire [6:0] _T_584 = _T_127 ? 7'h0 : _T_583; // @[Lookup.scala 33:37]
  wire [6:0] _T_585 = _T_125 ? 7'hf : _T_584; // @[Lookup.scala 33:37]
  wire [6:0] _T_586 = _T_123 ? 7'he : _T_585; // @[Lookup.scala 33:37]
  wire [6:0] _T_587 = _T_121 ? 7'hd : _T_586; // @[Lookup.scala 33:37]
  wire [6:0] _T_588 = _T_119 ? 7'hc : _T_587; // @[Lookup.scala 33:37]
  wire [6:0] _T_589 = _T_117 ? 7'h8 : _T_588; // @[Lookup.scala 33:37]
  wire [6:0] _T_590 = _T_115 ? 7'h7 : _T_589; // @[Lookup.scala 33:37]
  wire [6:0] _T_591 = _T_113 ? 7'h6 : _T_590; // @[Lookup.scala 33:37]
  wire [6:0] _T_592 = _T_111 ? 7'h5 : _T_591; // @[Lookup.scala 33:37]
  wire [6:0] _T_593 = _T_109 ? 7'h4 : _T_592; // @[Lookup.scala 33:37]
  wire [6:0] _T_594 = _T_107 ? 7'h3 : _T_593; // @[Lookup.scala 33:37]
  wire [6:0] _T_595 = _T_105 ? 7'h2 : _T_594; // @[Lookup.scala 33:37]
  wire [6:0] _T_596 = _T_103 ? 7'h1 : _T_595; // @[Lookup.scala 33:37]
  wire [6:0] _T_597 = _T_101 ? 7'h0 : _T_596; // @[Lookup.scala 33:37]
  wire [6:0] _T_598 = _T_99 ? 7'h2 : _T_597; // @[Lookup.scala 33:37]
  wire [6:0] _T_599 = _T_97 ? 7'hb : _T_598; // @[Lookup.scala 33:37]
  wire [6:0] _T_600 = _T_95 ? 7'h3 : _T_599; // @[Lookup.scala 33:37]
  wire [6:0] _T_601 = _T_93 ? 7'h6 : _T_600; // @[Lookup.scala 33:37]
  wire [6:0] _T_602 = _T_91 ? 7'h28 : _T_601; // @[Lookup.scala 33:37]
  wire [6:0] _T_603 = _T_89 ? 7'h60 : _T_602; // @[Lookup.scala 33:37]
  wire [6:0] _T_604 = _T_87 ? 7'h2d : _T_603; // @[Lookup.scala 33:37]
  wire [6:0] _T_605 = _T_85 ? 7'h25 : _T_604; // @[Lookup.scala 33:37]
  wire [6:0] _T_606 = _T_83 ? 7'h21 : _T_605; // @[Lookup.scala 33:37]
  wire [6:0] _T_607 = _T_81 ? 7'h2d : _T_606; // @[Lookup.scala 33:37]
  wire [6:0] _T_608 = _T_79 ? 7'h25 : _T_607; // @[Lookup.scala 33:37]
  wire [6:0] _T_609 = _T_77 ? 7'h21 : _T_608; // @[Lookup.scala 33:37]
  wire [6:0] _T_610 = _T_75 ? 7'h60 : _T_609; // @[Lookup.scala 33:37]
  wire [6:0] _T_611 = _T_73 ? 7'ha : _T_610; // @[Lookup.scala 33:37]
  wire [6:0] _T_612 = _T_71 ? 7'h9 : _T_611; // @[Lookup.scala 33:37]
  wire [6:0] _T_613 = _T_69 ? 7'h8 : _T_612; // @[Lookup.scala 33:37]
  wire [6:0] _T_614 = _T_67 ? 7'h5 : _T_613; // @[Lookup.scala 33:37]
  wire [6:0] _T_615 = _T_65 ? 7'h4 : _T_614; // @[Lookup.scala 33:37]
  wire [6:0] _T_616 = _T_63 ? 7'h2 : _T_615; // @[Lookup.scala 33:37]
  wire [6:0] _T_617 = _T_61 ? 7'h1 : _T_616; // @[Lookup.scala 33:37]
  wire [6:0] _T_618 = _T_59 ? 7'h0 : _T_617; // @[Lookup.scala 33:37]
  wire [6:0] _T_619 = _T_57 ? 7'h17 : _T_618; // @[Lookup.scala 33:37]
  wire [6:0] _T_620 = _T_55 ? 7'h16 : _T_619; // @[Lookup.scala 33:37]
  wire [6:0] _T_621 = _T_53 ? 7'h15 : _T_620; // @[Lookup.scala 33:37]
  wire [6:0] _T_622 = _T_51 ? 7'h14 : _T_621; // @[Lookup.scala 33:37]
  wire [6:0] _T_623 = _T_49 ? 7'h11 : _T_622; // @[Lookup.scala 33:37]
  wire [6:0] _T_624 = _T_47 ? 7'h10 : _T_623; // @[Lookup.scala 33:37]
  wire [6:0] _T_625 = _T_45 ? 7'h5a : _T_624; // @[Lookup.scala 33:37]
  wire [6:0] _T_626 = _T_43 ? 7'h58 : _T_625; // @[Lookup.scala 33:37]
  wire [6:0] _T_627 = _T_41 ? 7'h40 : _T_626; // @[Lookup.scala 33:37]
  wire [6:0] _T_628 = _T_39 ? 7'h40 : _T_627; // @[Lookup.scala 33:37]
  wire [6:0] _T_629 = _T_37 ? 7'hd : _T_628; // @[Lookup.scala 33:37]
  wire [6:0] _T_630 = _T_35 ? 7'h8 : _T_629; // @[Lookup.scala 33:37]
  wire [6:0] _T_631 = _T_33 ? 7'h7 : _T_630; // @[Lookup.scala 33:37]
  wire [6:0] _T_632 = _T_31 ? 7'h6 : _T_631; // @[Lookup.scala 33:37]
  wire [6:0] _T_633 = _T_29 ? 7'h5 : _T_632; // @[Lookup.scala 33:37]
  wire [6:0] _T_634 = _T_27 ? 7'h4 : _T_633; // @[Lookup.scala 33:37]
  wire [6:0] _T_635 = _T_25 ? 7'h3 : _T_634; // @[Lookup.scala 33:37]
  wire [6:0] _T_636 = _T_23 ? 7'h2 : _T_635; // @[Lookup.scala 33:37]
  wire [6:0] _T_637 = _T_21 ? 7'h1 : _T_636; // @[Lookup.scala 33:37]
  wire [6:0] _T_638 = _T_19 ? 7'h40 : _T_637; // @[Lookup.scala 33:37]
  wire [6:0] _T_639 = _T_17 ? 7'hd : _T_638; // @[Lookup.scala 33:37]
  wire [6:0] _T_640 = _T_15 ? 7'h7 : _T_639; // @[Lookup.scala 33:37]
  wire [6:0] _T_641 = _T_13 ? 7'h6 : _T_640; // @[Lookup.scala 33:37]
  wire [6:0] _T_642 = _T_11 ? 7'h5 : _T_641; // @[Lookup.scala 33:37]
  wire [6:0] _T_643 = _T_9 ? 7'h4 : _T_642; // @[Lookup.scala 33:37]
  wire [6:0] _T_644 = _T_7 ? 7'h3 : _T_643; // @[Lookup.scala 33:37]
  wire [6:0] _T_645 = _T_5 ? 7'h2 : _T_644; // @[Lookup.scala 33:37]
  wire [6:0] _T_646 = _T_3 ? 7'h1 : _T_645; // @[Lookup.scala 33:37]
  wire [6:0] decodeList_2 = _T_1 ? 7'h40 : _T_646; // @[Lookup.scala 33:37]
  wire  hasIntr = |intrVecIDU; // @[IDU.scala 186:22]
  wire [3:0] instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h0 : decodeList_0; // @[IDU.scala 38:75]
  wire [2:0] fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[IDU.scala 38:75]
  wire [6:0] fuOpType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[IDU.scala 38:75]
  wire  isRVC = io_in_bits_instr[1:0] != 2'h3; // @[IDU.scala 40:45]
  wire [4:0] _T_720 = _T_193 ? 5'h3 : 5'h10; // @[Lookup.scala 33:37]
  wire [4:0] _T_721 = _T_191 ? 5'h2 : _T_720; // @[Lookup.scala 33:37]
  wire [4:0] _T_722 = _T_189 ? 5'h10 : _T_721; // @[Lookup.scala 33:37]
  wire [4:0] _T_723 = _T_187 ? 5'h10 : _T_722; // @[Lookup.scala 33:37]
  wire [4:0] _T_724 = _T_185 ? 5'hf : _T_723; // @[Lookup.scala 33:37]
  wire [4:0] _T_725 = _T_183 ? 5'h10 : _T_724; // @[Lookup.scala 33:37]
  wire [4:0] _T_726 = _T_181 ? 5'h10 : _T_725; // @[Lookup.scala 33:37]
  wire [4:0] _T_727 = _T_179 ? 5'h1 : _T_726; // @[Lookup.scala 33:37]
  wire [4:0] _T_728 = _T_177 ? 5'h0 : _T_727; // @[Lookup.scala 33:37]
  wire [4:0] _T_729 = _T_175 ? 5'ha : _T_728; // @[Lookup.scala 33:37]
  wire [4:0] _T_730 = _T_173 ? 5'h9 : _T_729; // @[Lookup.scala 33:37]
  wire [4:0] _T_731 = _T_171 ? 5'h9 : _T_730; // @[Lookup.scala 33:37]
  wire [4:0] _T_732 = _T_169 ? 5'h8 : _T_731; // @[Lookup.scala 33:37]
  wire [4:0] _T_733 = _T_167 ? 5'h10 : _T_732; // @[Lookup.scala 33:37]
  wire [4:0] _T_734 = _T_165 ? 5'h10 : _T_733; // @[Lookup.scala 33:37]
  wire [4:0] _T_735 = _T_163 ? 5'h10 : _T_734; // @[Lookup.scala 33:37]
  wire [4:0] _T_736 = _T_161 ? 5'h10 : _T_735; // @[Lookup.scala 33:37]
  wire [4:0] _T_737 = _T_159 ? 5'h10 : _T_736; // @[Lookup.scala 33:37]
  wire [4:0] _T_738 = _T_157 ? 5'h10 : _T_737; // @[Lookup.scala 33:37]
  wire [4:0] _T_739 = _T_155 ? 5'ha : _T_738; // @[Lookup.scala 33:37]
  wire [4:0] _T_740 = _T_153 ? 5'ha : _T_739; // @[Lookup.scala 33:37]
  wire [4:0] _T_741 = _T_151 ? 5'ha : _T_740; // @[Lookup.scala 33:37]
  wire [4:0] _T_742 = _T_149 ? 5'hb : _T_741; // @[Lookup.scala 33:37]
  wire [4:0] _T_743 = _T_147 ? 5'hd : _T_742; // @[Lookup.scala 33:37]
  wire [4:0] _T_744 = _T_145 ? 5'ha : _T_743; // @[Lookup.scala 33:37]
  wire [4:0] _T_745 = _T_143 ? 5'hc : _T_744; // @[Lookup.scala 33:37]
  wire [4:0] _T_746 = _T_141 ? 5'hc : _T_745; // @[Lookup.scala 33:37]
  wire [4:0] _T_747 = _T_139 ? 5'h10 : _T_746; // @[Lookup.scala 33:37]
  wire [4:0] _T_748 = _T_137 ? 5'h5 : _T_747; // @[Lookup.scala 33:37]
  wire [4:0] _T_749 = _T_135 ? 5'h4 : _T_748; // @[Lookup.scala 33:37]
  wire [4:0] _T_750 = _T_133 ? 5'h7 : _T_749; // @[Lookup.scala 33:37]
  wire [4:0] _T_751 = _T_131 ? 5'h6 : _T_750; // @[Lookup.scala 33:37]
  wire [4:0] rvcImmType = _T_129 ? 5'he : _T_751; // @[Lookup.scala 33:37]
  wire [3:0] _T_752 = _T_193 ? 4'h9 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_753 = _T_191 ? 4'h9 : _T_752; // @[Lookup.scala 33:37]
  wire [3:0] _T_754 = _T_189 ? 4'h2 : _T_753; // @[Lookup.scala 33:37]
  wire [3:0] _T_755 = _T_187 ? 4'h4 : _T_754; // @[Lookup.scala 33:37]
  wire [3:0] _T_756 = _T_185 ? 4'h0 : _T_755; // @[Lookup.scala 33:37]
  wire [3:0] _T_757 = _T_183 ? 4'h5 : _T_756; // @[Lookup.scala 33:37]
  wire [3:0] _T_758 = _T_181 ? 4'h4 : _T_757; // @[Lookup.scala 33:37]
  wire [3:0] _T_759 = _T_179 ? 4'h9 : _T_758; // @[Lookup.scala 33:37]
  wire [3:0] _T_760 = _T_177 ? 4'h9 : _T_759; // @[Lookup.scala 33:37]
  wire [3:0] _T_761 = _T_175 ? 4'h2 : _T_760; // @[Lookup.scala 33:37]
  wire [3:0] _T_762 = _T_173 ? 4'h6 : _T_761; // @[Lookup.scala 33:37]
  wire [3:0] _T_763 = _T_171 ? 4'h6 : _T_762; // @[Lookup.scala 33:37]
  wire [3:0] _T_764 = _T_169 ? 4'h0 : _T_763; // @[Lookup.scala 33:37]
  wire [3:0] _T_765 = _T_167 ? 4'h6 : _T_764; // @[Lookup.scala 33:37]
  wire [3:0] _T_766 = _T_165 ? 4'h6 : _T_765; // @[Lookup.scala 33:37]
  wire [3:0] _T_767 = _T_163 ? 4'h6 : _T_766; // @[Lookup.scala 33:37]
  wire [3:0] _T_768 = _T_161 ? 4'h6 : _T_767; // @[Lookup.scala 33:37]
  wire [3:0] _T_769 = _T_159 ? 4'h6 : _T_768; // @[Lookup.scala 33:37]
  wire [3:0] _T_770 = _T_157 ? 4'h6 : _T_769; // @[Lookup.scala 33:37]
  wire [3:0] _T_771 = _T_155 ? 4'h6 : _T_770; // @[Lookup.scala 33:37]
  wire [3:0] _T_772 = _T_153 ? 4'h6 : _T_771; // @[Lookup.scala 33:37]
  wire [3:0] _T_773 = _T_151 ? 4'h6 : _T_772; // @[Lookup.scala 33:37]
  wire [3:0] _T_774 = _T_149 ? 4'h0 : _T_773; // @[Lookup.scala 33:37]
  wire [3:0] _T_775 = _T_147 ? 4'h9 : _T_774; // @[Lookup.scala 33:37]
  wire [3:0] _T_776 = _T_145 ? 4'h0 : _T_775; // @[Lookup.scala 33:37]
  wire [3:0] _T_777 = _T_143 ? 4'h2 : _T_776; // @[Lookup.scala 33:37]
  wire [3:0] _T_778 = _T_141 ? 4'h2 : _T_777; // @[Lookup.scala 33:37]
  wire [3:0] _T_779 = _T_139 ? 4'h0 : _T_778; // @[Lookup.scala 33:37]
  wire [3:0] _T_780 = _T_137 ? 4'h6 : _T_779; // @[Lookup.scala 33:37]
  wire [3:0] _T_781 = _T_135 ? 4'h6 : _T_780; // @[Lookup.scala 33:37]
  wire [3:0] _T_782 = _T_133 ? 4'h6 : _T_781; // @[Lookup.scala 33:37]
  wire [3:0] _T_783 = _T_131 ? 4'h6 : _T_782; // @[Lookup.scala 33:37]
  wire [3:0] rvcSrc1Type = _T_129 ? 4'h9 : _T_783; // @[Lookup.scala 33:37]
  wire [2:0] _T_784 = _T_193 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_785 = _T_191 ? 3'h5 : _T_784; // @[Lookup.scala 33:37]
  wire [2:0] _T_786 = _T_189 ? 3'h5 : _T_785; // @[Lookup.scala 33:37]
  wire [2:0] _T_787 = _T_187 ? 3'h0 : _T_786; // @[Lookup.scala 33:37]
  wire [2:0] _T_788 = _T_185 ? 3'h0 : _T_787; // @[Lookup.scala 33:37]
  wire [2:0] _T_789 = _T_183 ? 3'h0 : _T_788; // @[Lookup.scala 33:37]
  wire [2:0] _T_790 = _T_181 ? 3'h0 : _T_789; // @[Lookup.scala 33:37]
  wire [2:0] _T_791 = _T_179 ? 3'h0 : _T_790; // @[Lookup.scala 33:37]
  wire [2:0] _T_792 = _T_177 ? 3'h0 : _T_791; // @[Lookup.scala 33:37]
  wire [2:0] _T_793 = _T_175 ? 3'h0 : _T_792; // @[Lookup.scala 33:37]
  wire [2:0] _T_794 = _T_173 ? 3'h0 : _T_793; // @[Lookup.scala 33:37]
  wire [2:0] _T_795 = _T_171 ? 3'h0 : _T_794; // @[Lookup.scala 33:37]
  wire [2:0] _T_796 = _T_169 ? 3'h0 : _T_795; // @[Lookup.scala 33:37]
  wire [2:0] _T_797 = _T_167 ? 3'h7 : _T_796; // @[Lookup.scala 33:37]
  wire [2:0] _T_798 = _T_165 ? 3'h7 : _T_797; // @[Lookup.scala 33:37]
  wire [2:0] _T_799 = _T_163 ? 3'h7 : _T_798; // @[Lookup.scala 33:37]
  wire [2:0] _T_800 = _T_161 ? 3'h7 : _T_799; // @[Lookup.scala 33:37]
  wire [2:0] _T_801 = _T_159 ? 3'h7 : _T_800; // @[Lookup.scala 33:37]
  wire [2:0] _T_802 = _T_157 ? 3'h7 : _T_801; // @[Lookup.scala 33:37]
  wire [2:0] _T_803 = _T_155 ? 3'h0 : _T_802; // @[Lookup.scala 33:37]
  wire [2:0] _T_804 = _T_153 ? 3'h0 : _T_803; // @[Lookup.scala 33:37]
  wire [2:0] _T_805 = _T_151 ? 3'h0 : _T_804; // @[Lookup.scala 33:37]
  wire [2:0] _T_806 = _T_149 ? 3'h0 : _T_805; // @[Lookup.scala 33:37]
  wire [2:0] _T_807 = _T_147 ? 3'h0 : _T_806; // @[Lookup.scala 33:37]
  wire [2:0] _T_808 = _T_145 ? 3'h0 : _T_807; // @[Lookup.scala 33:37]
  wire [2:0] _T_809 = _T_143 ? 3'h0 : _T_808; // @[Lookup.scala 33:37]
  wire [2:0] _T_810 = _T_141 ? 3'h0 : _T_809; // @[Lookup.scala 33:37]
  wire [2:0] _T_811 = _T_139 ? 3'h0 : _T_810; // @[Lookup.scala 33:37]
  wire [2:0] _T_812 = _T_137 ? 3'h7 : _T_811; // @[Lookup.scala 33:37]
  wire [2:0] _T_813 = _T_135 ? 3'h7 : _T_812; // @[Lookup.scala 33:37]
  wire [2:0] _T_814 = _T_133 ? 3'h0 : _T_813; // @[Lookup.scala 33:37]
  wire [2:0] _T_815 = _T_131 ? 3'h0 : _T_814; // @[Lookup.scala 33:37]
  wire [2:0] rvcSrc2Type = _T_129 ? 3'h0 : _T_815; // @[Lookup.scala 33:37]
  wire [1:0] _T_818 = _T_189 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_819 = _T_187 ? 4'h8 : {{2'd0}, _T_818}; // @[Lookup.scala 33:37]
  wire [3:0] _T_820 = _T_185 ? 4'h0 : _T_819; // @[Lookup.scala 33:37]
  wire [3:0] _T_821 = _T_183 ? 4'h2 : _T_820; // @[Lookup.scala 33:37]
  wire [3:0] _T_822 = _T_181 ? 4'h0 : _T_821; // @[Lookup.scala 33:37]
  wire [3:0] _T_823 = _T_179 ? 4'h2 : _T_822; // @[Lookup.scala 33:37]
  wire [3:0] _T_824 = _T_177 ? 4'h2 : _T_823; // @[Lookup.scala 33:37]
  wire [3:0] _T_825 = _T_175 ? 4'h2 : _T_824; // @[Lookup.scala 33:37]
  wire [3:0] _T_826 = _T_173 ? 4'h0 : _T_825; // @[Lookup.scala 33:37]
  wire [3:0] _T_827 = _T_171 ? 4'h0 : _T_826; // @[Lookup.scala 33:37]
  wire [3:0] _T_828 = _T_169 ? 4'h0 : _T_827; // @[Lookup.scala 33:37]
  wire [3:0] _T_829 = _T_167 ? 4'h6 : _T_828; // @[Lookup.scala 33:37]
  wire [3:0] _T_830 = _T_165 ? 4'h6 : _T_829; // @[Lookup.scala 33:37]
  wire [3:0] _T_831 = _T_163 ? 4'h6 : _T_830; // @[Lookup.scala 33:37]
  wire [3:0] _T_832 = _T_161 ? 4'h6 : _T_831; // @[Lookup.scala 33:37]
  wire [3:0] _T_833 = _T_159 ? 4'h6 : _T_832; // @[Lookup.scala 33:37]
  wire [3:0] _T_834 = _T_157 ? 4'h6 : _T_833; // @[Lookup.scala 33:37]
  wire [3:0] _T_835 = _T_155 ? 4'h6 : _T_834; // @[Lookup.scala 33:37]
  wire [3:0] _T_836 = _T_153 ? 4'h6 : _T_835; // @[Lookup.scala 33:37]
  wire [3:0] _T_837 = _T_151 ? 4'h6 : _T_836; // @[Lookup.scala 33:37]
  wire [3:0] _T_838 = _T_149 ? 4'h2 : _T_837; // @[Lookup.scala 33:37]
  wire [3:0] _T_839 = _T_147 ? 4'h9 : _T_838; // @[Lookup.scala 33:37]
  wire [3:0] _T_840 = _T_145 ? 4'h2 : _T_839; // @[Lookup.scala 33:37]
  wire [3:0] _T_841 = _T_143 ? 4'h2 : _T_840; // @[Lookup.scala 33:37]
  wire [3:0] _T_842 = _T_141 ? 4'h2 : _T_841; // @[Lookup.scala 33:37]
  wire [3:0] _T_843 = _T_139 ? 4'h0 : _T_842; // @[Lookup.scala 33:37]
  wire [3:0] _T_844 = _T_137 ? 4'h0 : _T_843; // @[Lookup.scala 33:37]
  wire [3:0] _T_845 = _T_135 ? 4'h0 : _T_844; // @[Lookup.scala 33:37]
  wire [3:0] _T_846 = _T_133 ? 4'h7 : _T_845; // @[Lookup.scala 33:37]
  wire [3:0] _T_847 = _T_131 ? 4'h7 : _T_846; // @[Lookup.scala 33:37]
  wire [3:0] rvcDestType = _T_129 ? 4'h7 : _T_847; // @[Lookup.scala 33:37]
  wire  _T_848 = 4'h4 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_850 = 4'h2 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_851 = 4'hf == instrType; // @[LookupTree.scala 24:34]
  wire  _T_852 = 4'h1 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_853 = 4'h6 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_854 = 4'h7 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_855 = 4'h0 == instrType; // @[LookupTree.scala 24:34]
  wire  src1Type = _T_853 | _T_854 | _T_855; // @[Mux.scala 27:72]
  wire  src2Type = _T_848 | _T_853 | _T_854 | _T_855; // @[Mux.scala 27:72]
  wire [4:0] rs = io_in_bits_instr[19:15]; // @[IDU.scala 62:28]
  wire [4:0] rt = io_in_bits_instr[24:20]; // @[IDU.scala 62:43]
  wire [4:0] rd = io_in_bits_instr[11:7]; // @[IDU.scala 62:58]
  wire [4:0] rs2 = io_in_bits_instr[6:2]; // @[IDU.scala 65:24]
  wire  _T_895 = 3'h0 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_896 = 3'h1 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_897 = 3'h2 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_898 = 3'h3 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_899 = 3'h4 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_900 = 3'h5 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_901 = 3'h6 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_902 = 3'h7 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_903 = _T_895 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_904 = _T_896 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_905 = _T_897 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_906 = _T_898 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_907 = _T_899 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_908 = _T_900 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_909 = _T_901 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_910 = _T_902 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_911 = _T_903 | _T_904; // @[Mux.scala 27:72]
  wire [3:0] _T_912 = _T_911 | _T_905; // @[Mux.scala 27:72]
  wire [3:0] _T_913 = _T_912 | _T_906; // @[Mux.scala 27:72]
  wire [3:0] _T_914 = _T_913 | _T_907; // @[Mux.scala 27:72]
  wire [3:0] _T_915 = _T_914 | _T_908; // @[Mux.scala 27:72]
  wire [3:0] _T_916 = _T_915 | _T_909; // @[Mux.scala 27:72]
  wire [3:0] rs1p = _T_916 | _T_910; // @[Mux.scala 27:72]
  wire  _T_919 = 3'h0 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_920 = 3'h1 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_921 = 3'h2 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_922 = 3'h3 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_923 = 3'h4 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_924 = 3'h5 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_925 = 3'h6 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_926 = 3'h7 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_927 = _T_919 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_928 = _T_920 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_929 = _T_921 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_930 = _T_922 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_931 = _T_923 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_932 = _T_924 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_933 = _T_925 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_934 = _T_926 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_935 = _T_927 | _T_928; // @[Mux.scala 27:72]
  wire [3:0] _T_936 = _T_935 | _T_929; // @[Mux.scala 27:72]
  wire [3:0] _T_937 = _T_936 | _T_930; // @[Mux.scala 27:72]
  wire [3:0] _T_938 = _T_937 | _T_931; // @[Mux.scala 27:72]
  wire [3:0] _T_939 = _T_938 | _T_932; // @[Mux.scala 27:72]
  wire [3:0] _T_940 = _T_939 | _T_933; // @[Mux.scala 27:72]
  wire [3:0] rs2p = _T_940 | _T_934; // @[Mux.scala 27:72]
  wire [5:0] rvc_shamt = {io_in_bits_instr[12],rs2}; // @[Cat.scala 30:58]
  wire  _T_945 = 4'h3 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_946 = 4'h1 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_947 = 4'h2 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_948 = 4'h4 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_949 = 4'h5 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_950 = 4'h6 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_951 = 4'h7 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_952 = 4'h8 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_953 = 4'h9 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire [4:0] _T_955 = _T_945 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_956 = _T_946 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_957 = _T_947 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_958 = _T_948 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_959 = _T_949 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_960 = _T_950 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_961 = _T_951 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_963 = _T_953 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_965 = _T_955 | _T_956; // @[Mux.scala 27:72]
  wire [4:0] _T_966 = _T_965 | _T_957; // @[Mux.scala 27:72]
  wire [4:0] _T_967 = _T_966 | _T_958; // @[Mux.scala 27:72]
  wire [4:0] _T_968 = _T_967 | _T_959; // @[Mux.scala 27:72]
  wire [4:0] _GEN_9 = {{1'd0}, _T_960}; // @[Mux.scala 27:72]
  wire [4:0] _T_969 = _T_968 | _GEN_9; // @[Mux.scala 27:72]
  wire [4:0] _GEN_10 = {{1'd0}, _T_961}; // @[Mux.scala 27:72]
  wire [4:0] _T_970 = _T_969 | _GEN_10; // @[Mux.scala 27:72]
  wire [4:0] _GEN_11 = {{4'd0}, _T_952}; // @[Mux.scala 27:72]
  wire [4:0] _T_971 = _T_970 | _GEN_11; // @[Mux.scala 27:72]
  wire [4:0] _GEN_12 = {{3'd0}, _T_963}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src1 = _T_971 | _GEN_12; // @[Mux.scala 27:72]
  wire  _T_974 = 3'h3 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_975 = 3'h1 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_976 = 3'h2 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_977 = 3'h4 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_978 = 3'h5 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_979 = 3'h6 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_980 = 3'h7 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire [3:0] _GEN_13 = {{1'd0}, rvcSrc2Type}; // @[LookupTree.scala 24:34]
  wire  _T_981 = 4'h8 == _GEN_13; // @[LookupTree.scala 24:34]
  wire  _T_982 = 4'h9 == _GEN_13; // @[LookupTree.scala 24:34]
  wire [4:0] _T_984 = _T_974 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_985 = _T_975 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_986 = _T_976 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_987 = _T_977 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_988 = _T_978 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_989 = _T_979 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_990 = _T_980 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_992 = _T_982 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_994 = _T_984 | _T_985; // @[Mux.scala 27:72]
  wire [4:0] _T_995 = _T_994 | _T_986; // @[Mux.scala 27:72]
  wire [4:0] _T_996 = _T_995 | _T_987; // @[Mux.scala 27:72]
  wire [4:0] _T_997 = _T_996 | _T_988; // @[Mux.scala 27:72]
  wire [4:0] _GEN_15 = {{1'd0}, _T_989}; // @[Mux.scala 27:72]
  wire [4:0] _T_998 = _T_997 | _GEN_15; // @[Mux.scala 27:72]
  wire [4:0] _GEN_16 = {{1'd0}, _T_990}; // @[Mux.scala 27:72]
  wire [4:0] _T_999 = _T_998 | _GEN_16; // @[Mux.scala 27:72]
  wire [4:0] _GEN_17 = {{4'd0}, _T_981}; // @[Mux.scala 27:72]
  wire [4:0] _T_1000 = _T_999 | _GEN_17; // @[Mux.scala 27:72]
  wire [4:0] _GEN_18 = {{3'd0}, _T_992}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src2 = _T_1000 | _GEN_18; // @[Mux.scala 27:72]
  wire  _T_1003 = 4'h3 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1004 = 4'h1 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1005 = 4'h2 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1006 = 4'h4 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1007 = 4'h5 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1008 = 4'h6 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1009 = 4'h7 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1010 = 4'h8 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1011 = 4'h9 == rvcDestType; // @[LookupTree.scala 24:34]
  wire [4:0] _T_1013 = _T_1003 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1014 = _T_1004 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1015 = _T_1005 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1016 = _T_1006 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1017 = _T_1007 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1018 = _T_1008 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1019 = _T_1009 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_1021 = _T_1011 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1023 = _T_1013 | _T_1014; // @[Mux.scala 27:72]
  wire [4:0] _T_1024 = _T_1023 | _T_1015; // @[Mux.scala 27:72]
  wire [4:0] _T_1025 = _T_1024 | _T_1016; // @[Mux.scala 27:72]
  wire [4:0] _T_1026 = _T_1025 | _T_1017; // @[Mux.scala 27:72]
  wire [4:0] _GEN_19 = {{1'd0}, _T_1018}; // @[Mux.scala 27:72]
  wire [4:0] _T_1027 = _T_1026 | _GEN_19; // @[Mux.scala 27:72]
  wire [4:0] _GEN_20 = {{1'd0}, _T_1019}; // @[Mux.scala 27:72]
  wire [4:0] _T_1028 = _T_1027 | _GEN_20; // @[Mux.scala 27:72]
  wire [4:0] _GEN_21 = {{4'd0}, _T_1010}; // @[Mux.scala 27:72]
  wire [4:0] _T_1029 = _T_1028 | _GEN_21; // @[Mux.scala 27:72]
  wire [4:0] _GEN_22 = {{3'd0}, _T_1021}; // @[Mux.scala 27:72]
  wire [4:0] rvc_dest = _T_1029 | _GEN_22; // @[Mux.scala 27:72]
  wire [4:0] rfSrc1 = isRVC ? rvc_src1 : rs; // @[IDU.scala 89:19]
  wire [4:0] rfSrc2 = isRVC ? rvc_src2 : rt; // @[IDU.scala 90:19]
  wire [4:0] rfDest = isRVC ? rvc_dest : rd; // @[IDU.scala 91:19]
  wire [4:0] _T_1037 = instrType[2] ? rfDest : 5'h0; // @[IDU.scala 97:33]
  wire [51:0] _T_1041 = io_in_bits_instr[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1042 = {_T_1041,io_in_bits_instr[31:20]}; // @[Cat.scala 30:58]
  wire [11:0] _T_1045 = {io_in_bits_instr[31:25],rd}; // @[Cat.scala 30:58]
  wire [51:0] _T_1048 = _T_1045[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1049 = {_T_1048,io_in_bits_instr[31:25],rd}; // @[Cat.scala 30:58]
  wire [12:0] _T_1061 = {io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}; // @[Cat.scala 30:58]
  wire [50:0] _T_1064 = _T_1061[12] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1065 = {_T_1064,io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8]
    ,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_1067 = {io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_1070 = _T_1067[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1071 = {_T_1070,io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 30:58]
  wire [20:0] _T_1076 = {io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0}
    ; // @[Cat.scala 30:58]
  wire [42:0] _T_1079 = _T_1076[20] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1080 = {_T_1079,io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:
    21],1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1087 = _T_848 ? _T_1042 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1088 = _T_850 ? _T_1049 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1089 = _T_851 ? _T_1049 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1090 = _T_852 ? _T_1065 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1091 = _T_853 ? _T_1071 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1092 = _T_854 ? _T_1080 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1093 = _T_1087 | _T_1088; // @[Mux.scala 27:72]
  wire [63:0] _T_1094 = _T_1093 | _T_1089; // @[Mux.scala 27:72]
  wire [63:0] _T_1095 = _T_1094 | _T_1090; // @[Mux.scala 27:72]
  wire [63:0] _T_1096 = _T_1095 | _T_1091; // @[Mux.scala 27:72]
  wire [63:0] imm = _T_1096 | _T_1092; // @[Mux.scala 27:72]
  wire [63:0] _T_1102 = {56'h0,io_in_bits_instr[3:2],io_in_bits_instr[12],io_in_bits_instr[6:4],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1107 = {55'h0,io_in_bits_instr[4:2],io_in_bits_instr[12],io_in_bits_instr[6:5],3'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1111 = {56'h0,io_in_bits_instr[8:7],io_in_bits_instr[12:9],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1115 = {55'h0,io_in_bits_instr[9:7],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1120 = {57'h0,io_in_bits_instr[5],io_in_bits_instr[12:10],io_in_bits_instr[6],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1124 = {56'h0,io_in_bits_instr[6:5],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 30:58]
  wire [11:0] _T_1142 = {io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],
    io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 30:58]
  wire [51:0] _T_1145 = _T_1142[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1146 = {_T_1145,io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],
    io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 30:58]
  wire [8:0] _T_1152 = {io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],
    io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 30:58]
  wire [54:0] _T_1155 = _T_1152[8] ? 55'h7fffffffffffff : 55'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1156 = {_T_1155,io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],
    io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 30:58]
  wire [57:0] _T_1162 = rvc_shamt[5] ? 58'h3ffffffffffffff : 58'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1163 = {_T_1162,io_in_bits_instr[12],rs2}; // @[Cat.scala 30:58]
  wire [17:0] _T_1166 = {io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 30:58]
  wire [45:0] _T_1169 = _T_1166[17] ? 46'h3fffffffffff : 46'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1170 = {_T_1169,io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 30:58]
  wire [9:0] _T_1183 = {io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],
    io_in_bits_instr[6],4'h0}; // @[Cat.scala 30:58]
  wire [53:0] _T_1186 = _T_1183[9] ? 54'h3fffffffffffff : 54'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1187 = {_T_1186,io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],
    io_in_bits_instr[6],4'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1193 = {54'h0,io_in_bits_instr[10:7],io_in_bits_instr[12:11],io_in_bits_instr[5],io_in_bits_instr[6],2'h0
    }; // @[Cat.scala 30:58]
  wire  _T_1195 = 5'h0 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1196 = 5'h1 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1197 = 5'h2 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1198 = 5'h3 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1199 = 5'h4 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1200 = 5'h5 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1201 = 5'h6 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1202 = 5'h7 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1203 = 5'h8 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1204 = 5'h9 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1205 = 5'ha == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1206 = 5'hb == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1207 = 5'hc == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1208 = 5'hd == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1209 = 5'he == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1210 = 5'hf == rvcImmType; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1212 = _T_1195 ? _T_1102 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1213 = _T_1196 ? _T_1107 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1214 = _T_1197 ? _T_1111 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1215 = _T_1198 ? _T_1115 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1216 = _T_1199 ? _T_1120 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1217 = _T_1200 ? _T_1124 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1218 = _T_1201 ? _T_1120 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1219 = _T_1202 ? _T_1124 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1220 = _T_1203 ? _T_1146 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1221 = _T_1204 ? _T_1156 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1222 = _T_1205 ? _T_1163 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1223 = _T_1206 ? _T_1170 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1224 = _T_1207 ? _T_1163 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1225 = _T_1208 ? _T_1187 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1226 = _T_1209 ? _T_1193 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1227 = _T_1210 ? 64'h1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1229 = _T_1212 | _T_1213; // @[Mux.scala 27:72]
  wire [63:0] _T_1230 = _T_1229 | _T_1214; // @[Mux.scala 27:72]
  wire [63:0] _T_1231 = _T_1230 | _T_1215; // @[Mux.scala 27:72]
  wire [63:0] _T_1232 = _T_1231 | _T_1216; // @[Mux.scala 27:72]
  wire [63:0] _T_1233 = _T_1232 | _T_1217; // @[Mux.scala 27:72]
  wire [63:0] _T_1234 = _T_1233 | _T_1218; // @[Mux.scala 27:72]
  wire [63:0] _T_1235 = _T_1234 | _T_1219; // @[Mux.scala 27:72]
  wire [63:0] _T_1236 = _T_1235 | _T_1220; // @[Mux.scala 27:72]
  wire [63:0] _T_1237 = _T_1236 | _T_1221; // @[Mux.scala 27:72]
  wire [63:0] _T_1238 = _T_1237 | _T_1222; // @[Mux.scala 27:72]
  wire [63:0] _T_1239 = _T_1238 | _T_1223; // @[Mux.scala 27:72]
  wire [63:0] _T_1240 = _T_1239 | _T_1224; // @[Mux.scala 27:72]
  wire [63:0] _T_1241 = _T_1240 | _T_1225; // @[Mux.scala 27:72]
  wire [63:0] _T_1242 = _T_1241 | _T_1226; // @[Mux.scala 27:72]
  wire [63:0] immrvc = _T_1242 | _T_1227; // @[Mux.scala 27:72]
  wire  _T_1245 = fuType == 3'h0; // @[IDU.scala 132:16]
  wire  _T_1248 = rfDest == 5'h1 | rfDest == 5'h5; // @[IDU.scala 133:42]
  wire [6:0] _GEN_0 = _T_1248 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[IDU.scala 134:{57,85} 47:29]
  wire  _T_1254 = rfSrc1 == 5'h1 | rfSrc1 == 5'h5; // @[IDU.scala 133:42]
  wire [6:0] _GEN_1 = _T_1254 ? 7'h5e : _GEN_0; // @[IDU.scala 136:{29,57}]
  wire [6:0] _GEN_2 = _T_1248 ? 7'h5c : _GEN_1; // @[IDU.scala 137:{29,57}]
  wire [6:0] _GEN_3 = fuOpType == 7'h5a ? _GEN_2 : _GEN_0; // @[IDU.scala 135:40]
  wire  _T_1264 = ~io_in_bits_instr[14]; // @[IDU.scala 146:39]
  wire  _GEN_5 = _T_1264 ? 1'h0 : instrType[2]; // @[IDU.scala 148:27 149:32 96:27]
  wire [4:0] _GEN_6 = _T_1264 ? 5'h0 : _T_1037; // @[IDU.scala 148:27 150:32 97:27]
  wire  _T_1280 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_1281 = ~hasIntr; // @[IDU.scala 176:51]
  wire [7:0] _T_1319 = {7'h17 == fuOpType,7'h16 == fuOpType,7'h15 == fuOpType,7'h14 == fuOpType,7'h11 == fuOpType,7'h10
     == fuOpType,7'h5a == fuOpType,7'h58 == fuOpType}; // @[IDU.scala 202:84]
  assign io_in_ready = ~io_in_valid | _T_1280 & ~hasIntr; // @[IDU.scala 176:31]
  assign io_out_valid = io_in_valid; // @[IDU.scala 175:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[IDU.scala 177:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[IDU.scala 177:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[IDU.scala 177:18]
  assign io_out_bits_cf_exceptionVec_1 = |io_in_bits_pc[38:32] & ~DTLBENABLE; // @[IDU.scala 195:98]
  assign io_out_bits_cf_exceptionVec_2 = instrType == 4'h0 & _T_1281 & io_in_valid; // @[IDU.scala 192:83]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[IDU.scala 193:47]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[IDU.scala 185:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[IDU.scala 177:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_bits_crossPageIPFFix; // @[IDU.scala 177:18]
  assign io_out_bits_ctrl_src1Type = io_in_bits_instr[6:0] == 7'h37 ? 1'h0 : src1Type; // @[IDU.scala 141:35]
  assign io_out_bits_ctrl_src2Type = _T_848 | _T_853 | _T_854 | _T_855; // @[Mux.scala 27:72]
  assign io_out_bits_ctrl_fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 :
    decodeList_1; // @[IDU.scala 38:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 3'h0 ? _GEN_3 : fuOpType; // @[IDU.scala 132:32 47:29]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rfSrc1; // @[IDU.scala 94:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rfSrc2 : 5'h0; // @[IDU.scala 95:33]
  assign io_out_bits_ctrl_rfWen = fuType == 3'h5 ? _GEN_5 : instrType[2]; // @[IDU.scala 145:32 96:27]
  assign io_out_bits_ctrl_rfDest = fuType == 3'h5 ? _GEN_6 : _T_1037; // @[IDU.scala 145:32 97:27]
  assign io_out_bits_ctrl_vtag = io_in_bits_instr[26:24]; // @[IDU.scala 153:38]
  assign io_out_bits_ctrl_vec_addr = io_in_bits_instr[11:7]; // @[IDU.scala 154:38]
  assign io_out_bits_ctrl_length_k = io_in_bits_instr[23:20]; // @[IDU.scala 155:38]
  assign io_out_bits_ctrl_algorithm = io_in_bits_instr[16:15]; // @[IDU.scala 156:38]
  assign io_out_bits_data_imm = isRVC ? immrvc : imm; // @[IDU.scala 130:31]
  assign io_isBranch = |_T_1319 & _T_1245; // @[IDU.scala 202:95]
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_instr,
  input  [38:0] io_in_0_bits_pc,
  input  [38:0] io_in_0_bits_pnpc,
  input         io_in_0_bits_exceptionVec_12,
  input  [3:0]  io_in_0_bits_brIdx,
  input         io_in_0_bits_crossPageIPFFix,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output [63:0] io_out_0_bits_cf_runahead_checkpoint_id,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output [2:0]  io_out_0_bits_ctrl_vtag,
  output [4:0]  io_out_0_bits_ctrl_vec_addr,
  output [3:0]  io_out_0_bits_ctrl_length_k,
  output [1:0]  io_out_0_bits_ctrl_algorithm,
  output [63:0] io_out_0_bits_data_imm,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [63:0] io_out_1_bits_cf_instr,
  output [38:0] io_out_1_bits_cf_pc,
  output [38:0] io_out_1_bits_cf_pnpc,
  output        io_out_1_bits_cf_exceptionVec_1,
  output        io_out_1_bits_cf_exceptionVec_2,
  output        io_out_1_bits_cf_exceptionVec_12,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  output [3:0]  io_out_1_bits_cf_brIdx,
  output        io_out_1_bits_cf_crossPageIPFFix,
  output        io_out_1_bits_ctrl_src1Type,
  output        io_out_1_bits_ctrl_src2Type,
  output [2:0]  io_out_1_bits_ctrl_fuType,
  output [6:0]  io_out_1_bits_ctrl_fuOpType,
  output [4:0]  io_out_1_bits_ctrl_rfSrc1,
  output [4:0]  io_out_1_bits_ctrl_rfSrc2,
  output        io_out_1_bits_ctrl_rfWen,
  output [4:0]  io_out_1_bits_ctrl_rfDest,
  output [2:0]  io_out_1_bits_ctrl_vtag,
  output [4:0]  io_out_1_bits_ctrl_vec_addr,
  output [3:0]  io_out_1_bits_ctrl_length_k,
  output [1:0]  io_out_1_bits_ctrl_algorithm,
  output [63:0] io_out_1_bits_data_imm,
  input         vmEnable,
  input  [11:0] intrVec
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  decoder1_io_in_ready; // @[IDU.scala 211:25]
  wire  decoder1_io_in_valid; // @[IDU.scala 211:25]
  wire [63:0] decoder1_io_in_bits_instr; // @[IDU.scala 211:25]
  wire [38:0] decoder1_io_in_bits_pc; // @[IDU.scala 211:25]
  wire [38:0] decoder1_io_in_bits_pnpc; // @[IDU.scala 211:25]
  wire  decoder1_io_in_bits_exceptionVec_12; // @[IDU.scala 211:25]
  wire [3:0] decoder1_io_in_bits_brIdx; // @[IDU.scala 211:25]
  wire  decoder1_io_in_bits_crossPageIPFFix; // @[IDU.scala 211:25]
  wire  decoder1_io_out_ready; // @[IDU.scala 211:25]
  wire  decoder1_io_out_valid; // @[IDU.scala 211:25]
  wire [63:0] decoder1_io_out_bits_cf_instr; // @[IDU.scala 211:25]
  wire [38:0] decoder1_io_out_bits_cf_pc; // @[IDU.scala 211:25]
  wire [38:0] decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 211:25]
  wire [3:0] decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 211:25]
  wire [2:0] decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 211:25]
  wire [6:0] decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 211:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 211:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 211:25]
  wire  decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 211:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 211:25]
  wire [2:0] decoder1_io_out_bits_ctrl_vtag; // @[IDU.scala 211:25]
  wire [4:0] decoder1_io_out_bits_ctrl_vec_addr; // @[IDU.scala 211:25]
  wire [3:0] decoder1_io_out_bits_ctrl_length_k; // @[IDU.scala 211:25]
  wire [1:0] decoder1_io_out_bits_ctrl_algorithm; // @[IDU.scala 211:25]
  wire [63:0] decoder1_io_out_bits_data_imm; // @[IDU.scala 211:25]
  wire  decoder1_io_isBranch; // @[IDU.scala 211:25]
  wire  decoder1_DTLBENABLE; // @[IDU.scala 211:25]
  wire [11:0] decoder1_intrVecIDU; // @[IDU.scala 211:25]
  wire  decoder2_io_in_ready; // @[IDU.scala 212:25]
  wire  decoder2_io_in_valid; // @[IDU.scala 212:25]
  wire [63:0] decoder2_io_in_bits_instr; // @[IDU.scala 212:25]
  wire [38:0] decoder2_io_in_bits_pc; // @[IDU.scala 212:25]
  wire [38:0] decoder2_io_in_bits_pnpc; // @[IDU.scala 212:25]
  wire  decoder2_io_in_bits_exceptionVec_12; // @[IDU.scala 212:25]
  wire [3:0] decoder2_io_in_bits_brIdx; // @[IDU.scala 212:25]
  wire  decoder2_io_in_bits_crossPageIPFFix; // @[IDU.scala 212:25]
  wire  decoder2_io_out_ready; // @[IDU.scala 212:25]
  wire  decoder2_io_out_valid; // @[IDU.scala 212:25]
  wire [63:0] decoder2_io_out_bits_cf_instr; // @[IDU.scala 212:25]
  wire [38:0] decoder2_io_out_bits_cf_pc; // @[IDU.scala 212:25]
  wire [38:0] decoder2_io_out_bits_cf_pnpc; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 212:25]
  wire [3:0] decoder2_io_out_bits_cf_brIdx; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_ctrl_src1Type; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_ctrl_src2Type; // @[IDU.scala 212:25]
  wire [2:0] decoder2_io_out_bits_ctrl_fuType; // @[IDU.scala 212:25]
  wire [6:0] decoder2_io_out_bits_ctrl_fuOpType; // @[IDU.scala 212:25]
  wire [4:0] decoder2_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 212:25]
  wire [4:0] decoder2_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 212:25]
  wire  decoder2_io_out_bits_ctrl_rfWen; // @[IDU.scala 212:25]
  wire [4:0] decoder2_io_out_bits_ctrl_rfDest; // @[IDU.scala 212:25]
  wire [2:0] decoder2_io_out_bits_ctrl_vtag; // @[IDU.scala 212:25]
  wire [4:0] decoder2_io_out_bits_ctrl_vec_addr; // @[IDU.scala 212:25]
  wire [3:0] decoder2_io_out_bits_ctrl_length_k; // @[IDU.scala 212:25]
  wire [1:0] decoder2_io_out_bits_ctrl_algorithm; // @[IDU.scala 212:25]
  wire [63:0] decoder2_io_out_bits_data_imm; // @[IDU.scala 212:25]
  wire  decoder2_io_isBranch; // @[IDU.scala 212:25]
  wire  decoder2_DTLBENABLE; // @[IDU.scala 212:25]
  wire [11:0] decoder2_intrVecIDU; // @[IDU.scala 212:25]
  wire  runahead_io_clock; // @[IDU.scala 225:24]
  wire [7:0] runahead_io_coreid; // @[IDU.scala 225:24]
  wire [7:0] runahead_io_index; // @[IDU.scala 225:24]
  wire  runahead_io_valid; // @[IDU.scala 225:24]
  wire  runahead_io_branch; // @[IDU.scala 225:24]
  wire  runahead_io_may_replay; // @[IDU.scala 225:24]
  wire [63:0] runahead_io_pc; // @[IDU.scala 225:24]
  wire [63:0] runahead_io_checkpoint_id; // @[IDU.scala 225:24]
  reg [63:0] checkpoint_id; // @[IDU.scala 222:30]
  wire [63:0] _T_3 = checkpoint_id + 64'h1; // @[IDU.scala 233:36]
  Decoder decoder1 ( // @[IDU.scala 211:25]
    .io_in_ready(decoder1_io_in_ready),
    .io_in_valid(decoder1_io_in_valid),
    .io_in_bits_instr(decoder1_io_in_bits_instr),
    .io_in_bits_pc(decoder1_io_in_bits_pc),
    .io_in_bits_pnpc(decoder1_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder1_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder1_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder1_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder1_io_out_ready),
    .io_out_valid(decoder1_io_out_valid),
    .io_out_bits_cf_instr(decoder1_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder1_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder1_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder1_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder1_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder1_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder1_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder1_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder1_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder1_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder1_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder1_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder1_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder1_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder1_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder1_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder1_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder1_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder1_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder1_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_src1Type(decoder1_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder1_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder1_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder1_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder1_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder1_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder1_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder1_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_vtag(decoder1_io_out_bits_ctrl_vtag),
    .io_out_bits_ctrl_vec_addr(decoder1_io_out_bits_ctrl_vec_addr),
    .io_out_bits_ctrl_length_k(decoder1_io_out_bits_ctrl_length_k),
    .io_out_bits_ctrl_algorithm(decoder1_io_out_bits_ctrl_algorithm),
    .io_out_bits_data_imm(decoder1_io_out_bits_data_imm),
    .io_isBranch(decoder1_io_isBranch),
    .DTLBENABLE(decoder1_DTLBENABLE),
    .intrVecIDU(decoder1_intrVecIDU)
  );
  Decoder decoder2 ( // @[IDU.scala 212:25]
    .io_in_ready(decoder2_io_in_ready),
    .io_in_valid(decoder2_io_in_valid),
    .io_in_bits_instr(decoder2_io_in_bits_instr),
    .io_in_bits_pc(decoder2_io_in_bits_pc),
    .io_in_bits_pnpc(decoder2_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder2_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder2_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder2_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder2_io_out_ready),
    .io_out_valid(decoder2_io_out_valid),
    .io_out_bits_cf_instr(decoder2_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder2_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder2_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder2_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder2_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder2_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder2_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder2_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder2_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder2_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder2_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder2_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder2_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder2_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder2_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder2_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder2_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder2_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder2_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder2_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_src1Type(decoder2_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder2_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder2_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder2_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder2_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder2_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder2_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder2_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_vtag(decoder2_io_out_bits_ctrl_vtag),
    .io_out_bits_ctrl_vec_addr(decoder2_io_out_bits_ctrl_vec_addr),
    .io_out_bits_ctrl_length_k(decoder2_io_out_bits_ctrl_length_k),
    .io_out_bits_ctrl_algorithm(decoder2_io_out_bits_ctrl_algorithm),
    .io_out_bits_data_imm(decoder2_io_out_bits_data_imm),
    .io_isBranch(decoder2_io_isBranch),
    .DTLBENABLE(decoder2_DTLBENABLE),
    .intrVecIDU(decoder2_intrVecIDU)
  );
  DifftestRunaheadEvent runahead ( // @[IDU.scala 225:24]
    .io_clock(runahead_io_clock),
    .io_coreid(runahead_io_coreid),
    .io_index(runahead_io_index),
    .io_valid(runahead_io_valid),
    .io_branch(runahead_io_branch),
    .io_may_replay(runahead_io_may_replay),
    .io_pc(runahead_io_pc),
    .io_checkpoint_id(runahead_io_checkpoint_id)
  );
  assign io_in_0_ready = decoder1_io_in_ready; // @[IDU.scala 213:12]
  assign io_out_0_valid = decoder1_io_out_valid; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_instr = decoder1_io_out_bits_cf_instr; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_pc = decoder1_io_out_bits_cf_pc; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_pnpc = decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_0 = decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_2 = decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_4 = decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_6 = decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_8 = decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_10 = decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_brIdx = decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_crossPageIPFFix = decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 215:13]
  assign io_out_0_bits_cf_runahead_checkpoint_id = checkpoint_id; // @[IDU.scala 236:44]
  assign io_out_0_bits_ctrl_src1Type = decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_src2Type = decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_fuType = decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_rfWen = decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_rfDest = decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_vtag = decoder1_io_out_bits_ctrl_vtag; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_vec_addr = decoder1_io_out_bits_ctrl_vec_addr; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_length_k = decoder1_io_out_bits_ctrl_length_k; // @[IDU.scala 215:13]
  assign io_out_0_bits_ctrl_algorithm = decoder1_io_out_bits_ctrl_algorithm; // @[IDU.scala 215:13]
  assign io_out_0_bits_data_imm = decoder1_io_out_bits_data_imm; // @[IDU.scala 215:13]
  assign io_out_1_valid = decoder2_io_out_valid; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_instr = decoder2_io_out_bits_cf_instr; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_pc = decoder2_io_out_bits_cf_pc; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_pnpc = decoder2_io_out_bits_cf_pnpc; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_exceptionVec_1 = decoder2_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_exceptionVec_2 = decoder2_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_exceptionVec_12 = decoder2_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_0 = decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_1 = decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_2 = decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_3 = decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_4 = decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_5 = decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_6 = decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_7 = decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_8 = decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_9 = decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_10 = decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_intrVec_11 = decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_brIdx = decoder2_io_out_bits_cf_brIdx; // @[IDU.scala 216:13]
  assign io_out_1_bits_cf_crossPageIPFFix = decoder2_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_src1Type = decoder2_io_out_bits_ctrl_src1Type; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_src2Type = decoder2_io_out_bits_ctrl_src2Type; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_fuType = decoder2_io_out_bits_ctrl_fuType; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_fuOpType = decoder2_io_out_bits_ctrl_fuOpType; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_rfSrc1 = decoder2_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_rfSrc2 = decoder2_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_rfWen = decoder2_io_out_bits_ctrl_rfWen; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_rfDest = decoder2_io_out_bits_ctrl_rfDest; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_vtag = decoder2_io_out_bits_ctrl_vtag; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_vec_addr = decoder2_io_out_bits_ctrl_vec_addr; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_length_k = decoder2_io_out_bits_ctrl_length_k; // @[IDU.scala 216:13]
  assign io_out_1_bits_ctrl_algorithm = decoder2_io_out_bits_ctrl_algorithm; // @[IDU.scala 216:13]
  assign io_out_1_bits_data_imm = decoder2_io_out_bits_data_imm; // @[IDU.scala 216:13]
  assign decoder1_io_in_valid = io_in_0_valid; // @[IDU.scala 213:12]
  assign decoder1_io_in_bits_instr = io_in_0_bits_instr; // @[IDU.scala 213:12]
  assign decoder1_io_in_bits_pc = io_in_0_bits_pc; // @[IDU.scala 213:12]
  assign decoder1_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[IDU.scala 213:12]
  assign decoder1_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[IDU.scala 213:12]
  assign decoder1_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[IDU.scala 213:12]
  assign decoder1_io_in_bits_crossPageIPFFix = io_in_0_bits_crossPageIPFFix; // @[IDU.scala 213:12]
  assign decoder1_io_out_ready = io_out_0_ready; // @[IDU.scala 215:13]
  assign decoder1_DTLBENABLE = vmEnable;
  assign decoder1_intrVecIDU = intrVec;
  assign decoder2_io_in_valid = 1'h0; // @[IDU.scala 219:26]
  assign decoder2_io_in_bits_instr = 64'h0; // @[IDU.scala 214:12]
  assign decoder2_io_in_bits_pc = 39'h0; // @[IDU.scala 214:12]
  assign decoder2_io_in_bits_pnpc = 39'h0; // @[IDU.scala 214:12]
  assign decoder2_io_in_bits_exceptionVec_12 = 1'h0; // @[IDU.scala 214:12]
  assign decoder2_io_in_bits_brIdx = 4'h0; // @[IDU.scala 214:12]
  assign decoder2_io_in_bits_crossPageIPFFix = 1'h0; // @[IDU.scala 214:12]
  assign decoder2_io_out_ready = io_out_1_ready; // @[IDU.scala 216:13]
  assign decoder2_DTLBENABLE = vmEnable;
  assign decoder2_intrVecIDU = intrVec;
  assign runahead_io_clock = clock; // @[IDU.scala 226:29]
  assign runahead_io_coreid = 8'h0; // @[IDU.scala 227:29]
  assign runahead_io_index = 8'h0;
  assign runahead_io_valid = io_out_0_ready & io_out_0_valid; // @[Decoupled.scala 40:37]
  assign runahead_io_branch = decoder1_io_isBranch; // @[IDU.scala 229:29]
  assign runahead_io_may_replay = 1'h0;
  assign runahead_io_pc = {{25'd0}, io_out_0_bits_cf_pc}; // @[IDU.scala 230:29]
  assign runahead_io_checkpoint_id = checkpoint_id; // @[IDU.scala 231:29]
  always @(posedge clock) begin
    if (reset) begin // @[IDU.scala 222:30]
      checkpoint_id <= 64'h0; // @[IDU.scala 222:30]
    end else if (runahead_io_valid & runahead_io_branch) begin // @[IDU.scala 232:49]
      checkpoint_id <= _T_3; // @[IDU.scala 233:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  checkpoint_id = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_instr,
  input  [38:0] io_enq_bits_pc,
  input  [38:0] io_enq_bits_pnpc,
  input         io_enq_bits_exceptionVec_12,
  input  [3:0]  io_enq_bits_brIdx,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_instr,
  output [38:0] io_deq_bits_pc,
  output [38:0] io_deq_bits_pnpc,
  output        io_deq_bits_exceptionVec_12,
  output [3:0]  io_deq_bits_brIdx,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] MEM_instr [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_instr_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_instr_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [63:0] MEM_instr_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [63:0] MEM_instr_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_instr_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_instr_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_instr_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [38:0] MEM_pc [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_pc_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pc_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pc_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pc_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pc_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_pc_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_pc_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [38:0] MEM_pnpc [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_pnpc_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pnpc_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pnpc_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [38:0] MEM_pnpc_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_pnpc_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_pnpc_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_pnpc_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg  MEM_exceptionVec_12 [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_exceptionVec_12_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_exceptionVec_12_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_exceptionVec_12_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [3:0] MEM_brIdx [0:3]; // @[FlushableQueue.scala 23:24]
  wire  MEM_brIdx_MPORT_1_en; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_brIdx_MPORT_1_addr; // @[FlushableQueue.scala 23:24]
  wire [3:0] MEM_brIdx_MPORT_1_data; // @[FlushableQueue.scala 23:24]
  wire [3:0] MEM_brIdx_MPORT_data; // @[FlushableQueue.scala 23:24]
  wire [1:0] MEM_brIdx_MPORT_addr; // @[FlushableQueue.scala 23:24]
  wire  MEM_brIdx_MPORT_mask; // @[FlushableQueue.scala 23:24]
  wire  MEM_brIdx_MPORT_en; // @[FlushableQueue.scala 23:24]
  reg [1:0] value; // @[Counter.scala 60:40]
  reg [1:0] value_1; // @[Counter.scala 60:40]
  reg  REG; // @[FlushableQueue.scala 26:35]
  wire  _T = value == value_1; // @[FlushableQueue.scala 28:41]
  wire  _T_2 = _T & ~REG; // @[FlushableQueue.scala 29:33]
  wire  _T_3 = _T & REG; // @[FlushableQueue.scala 30:32]
  wire  _T_4 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _value_T_1 = value + 2'h1; // @[Counter.scala 76:24]
  wire [1:0] _value_T_3 = value_1 + 2'h1; // @[Counter.scala 76:24]
  assign MEM_instr_MPORT_1_en = 1'h1;
  assign MEM_instr_MPORT_1_addr = value_1;
  assign MEM_instr_MPORT_1_data = MEM_instr[MEM_instr_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_instr_MPORT_data = io_enq_bits_instr;
  assign MEM_instr_MPORT_addr = value;
  assign MEM_instr_MPORT_mask = 1'h1;
  assign MEM_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_pc_MPORT_1_en = 1'h1;
  assign MEM_pc_MPORT_1_addr = value_1;
  assign MEM_pc_MPORT_1_data = MEM_pc[MEM_pc_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_pc_MPORT_data = io_enq_bits_pc;
  assign MEM_pc_MPORT_addr = value;
  assign MEM_pc_MPORT_mask = 1'h1;
  assign MEM_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_pnpc_MPORT_1_en = 1'h1;
  assign MEM_pnpc_MPORT_1_addr = value_1;
  assign MEM_pnpc_MPORT_1_data = MEM_pnpc[MEM_pnpc_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_pnpc_MPORT_data = io_enq_bits_pnpc;
  assign MEM_pnpc_MPORT_addr = value;
  assign MEM_pnpc_MPORT_mask = 1'h1;
  assign MEM_pnpc_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_exceptionVec_12_MPORT_1_en = 1'h1;
  assign MEM_exceptionVec_12_MPORT_1_addr = value_1;
  assign MEM_exceptionVec_12_MPORT_1_data = MEM_exceptionVec_12[MEM_exceptionVec_12_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_exceptionVec_12_MPORT_data = io_enq_bits_exceptionVec_12;
  assign MEM_exceptionVec_12_MPORT_addr = value;
  assign MEM_exceptionVec_12_MPORT_mask = 1'h1;
  assign MEM_exceptionVec_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign MEM_brIdx_MPORT_1_en = 1'h1;
  assign MEM_brIdx_MPORT_1_addr = value_1;
  assign MEM_brIdx_MPORT_1_data = MEM_brIdx[MEM_brIdx_MPORT_1_addr]; // @[FlushableQueue.scala 23:24]
  assign MEM_brIdx_MPORT_data = io_enq_bits_brIdx;
  assign MEM_brIdx_MPORT_addr = value;
  assign MEM_brIdx_MPORT_mask = 1'h1;
  assign MEM_brIdx_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_3; // @[FlushableQueue.scala 46:19]
  assign io_deq_valid = ~_T_2; // @[FlushableQueue.scala 45:19]
  assign io_deq_bits_instr = MEM_instr_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_pc = MEM_pc_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_pnpc = MEM_pnpc_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_12 = MEM_exceptionVec_12_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  assign io_deq_bits_brIdx = MEM_brIdx_MPORT_1_data; // @[FlushableQueue.scala 47:15]
  always @(posedge clock) begin
    if (MEM_instr_MPORT_en & MEM_instr_MPORT_mask) begin
      MEM_instr[MEM_instr_MPORT_addr] <= MEM_instr_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_pc_MPORT_en & MEM_pc_MPORT_mask) begin
      MEM_pc[MEM_pc_MPORT_addr] <= MEM_pc_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_pnpc_MPORT_en & MEM_pnpc_MPORT_mask) begin
      MEM_pnpc[MEM_pnpc_MPORT_addr] <= MEM_pnpc_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_exceptionVec_12_MPORT_en & MEM_exceptionVec_12_MPORT_mask) begin
      MEM_exceptionVec_12[MEM_exceptionVec_12_MPORT_addr] <= MEM_exceptionVec_12_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (MEM_brIdx_MPORT_en & MEM_brIdx_MPORT_mask) begin
      MEM_brIdx[MEM_brIdx_MPORT_addr] <= MEM_brIdx_MPORT_data; // @[FlushableQueue.scala 23:24]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 2'h0; // @[Counter.scala 60:40]
    end else if (io_flush) begin // @[FlushableQueue.scala 62:19]
      value <= 2'h0; // @[FlushableQueue.scala 64:21]
    end else if (_T_4) begin // @[FlushableQueue.scala 34:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 2'h0; // @[Counter.scala 60:40]
    end else if (io_flush) begin // @[FlushableQueue.scala 62:19]
      value_1 <= 2'h0; // @[FlushableQueue.scala 65:21]
    end else if (_T_5) begin // @[FlushableQueue.scala 38:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[FlushableQueue.scala 26:35]
      REG <= 1'h0; // @[FlushableQueue.scala 26:35]
    end else if (io_flush) begin // @[FlushableQueue.scala 62:19]
      REG <= 1'h0; // @[FlushableQueue.scala 67:16]
    end else if (_T_4 != _T_5) begin // @[FlushableQueue.scala 41:28]
      REG <= _T_4; // @[FlushableQueue.scala 42:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_exceptionVec_12[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    MEM_brIdx[initvar] = _RAND_4[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  REG = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [86:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [86:0] io_imem_resp_bits_user,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output [63:0] io_out_0_bits_cf_runahead_checkpoint_id,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output [2:0]  io_out_0_bits_ctrl_vtag,
  output [4:0]  io_out_0_bits_ctrl_vec_addr,
  output [3:0]  io_out_0_bits_ctrl_length_k,
  output [1:0]  io_out_0_bits_ctrl_algorithm,
  output [63:0] io_out_0_bits_data_imm,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [63:0] io_out_1_bits_cf_instr,
  output [38:0] io_out_1_bits_cf_pc,
  output [38:0] io_out_1_bits_cf_pnpc,
  output        io_out_1_bits_cf_exceptionVec_1,
  output        io_out_1_bits_cf_exceptionVec_2,
  output        io_out_1_bits_cf_exceptionVec_12,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  output [3:0]  io_out_1_bits_cf_brIdx,
  output        io_out_1_bits_cf_crossPageIPFFix,
  output        io_out_1_bits_ctrl_src1Type,
  output        io_out_1_bits_ctrl_src2Type,
  output [2:0]  io_out_1_bits_ctrl_fuType,
  output [6:0]  io_out_1_bits_ctrl_fuOpType,
  output [4:0]  io_out_1_bits_ctrl_rfSrc1,
  output [4:0]  io_out_1_bits_ctrl_rfSrc2,
  output        io_out_1_bits_ctrl_rfWen,
  output [4:0]  io_out_1_bits_ctrl_rfDest,
  output [2:0]  io_out_1_bits_ctrl_vtag,
  output [4:0]  io_out_1_bits_ctrl_vec_addr,
  output [3:0]  io_out_1_bits_ctrl_length_k,
  output [1:0]  io_out_1_bits_ctrl_algorithm,
  output [63:0] io_out_1_bits_data_imm,
  output [3:0]  io_flushVec,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  input         io_ipf,
  input         flushICache,
  input         REG_0_valid,
  input  [38:0] REG_0_pc,
  input         REG_0_isMissPredict,
  input  [38:0] REG_0_actualTarget,
  input         REG_0_actualTaken,
  input  [6:0]  REG_0_fuOpType,
  input  [1:0]  REG_0_btbType,
  input         REG_0_isRVC,
  input         vmEnable,
  input  [11:0] intrVec,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[Frontend.scala 96:20]
  wire  ifu_reset; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_req_ready; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_req_valid; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[Frontend.scala 96:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_resp_ready; // @[Frontend.scala 96:20]
  wire  ifu_io_imem_resp_valid; // @[Frontend.scala 96:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[Frontend.scala 96:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[Frontend.scala 96:20]
  wire  ifu_io_out_ready; // @[Frontend.scala 96:20]
  wire  ifu_io_out_valid; // @[Frontend.scala 96:20]
  wire [63:0] ifu_io_out_bits_instr; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_out_bits_pc; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[Frontend.scala 96:20]
  wire  ifu_io_out_bits_exceptionVec_12; // @[Frontend.scala 96:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[Frontend.scala 96:20]
  wire [38:0] ifu_io_redirect_target; // @[Frontend.scala 96:20]
  wire  ifu_io_redirect_valid; // @[Frontend.scala 96:20]
  wire [3:0] ifu_io_flushVec; // @[Frontend.scala 96:20]
  wire  ifu_io_ipf; // @[Frontend.scala 96:20]
  wire  ifu_flushICache; // @[Frontend.scala 96:20]
  wire  ifu_REG_0_valid; // @[Frontend.scala 96:20]
  wire [38:0] ifu_REG_0_pc; // @[Frontend.scala 96:20]
  wire  ifu_REG_0_isMissPredict; // @[Frontend.scala 96:20]
  wire [38:0] ifu_REG_0_actualTarget; // @[Frontend.scala 96:20]
  wire  ifu_REG_0_actualTaken; // @[Frontend.scala 96:20]
  wire [6:0] ifu_REG_0_fuOpType; // @[Frontend.scala 96:20]
  wire [1:0] ifu_REG_0_btbType; // @[Frontend.scala 96:20]
  wire  ifu_REG_0_isRVC; // @[Frontend.scala 96:20]
  wire  ifu_flushTLB; // @[Frontend.scala 96:20]
  wire  ibf_clock; // @[Frontend.scala 97:19]
  wire  ibf_reset; // @[Frontend.scala 97:19]
  wire  ibf_io_in_ready; // @[Frontend.scala 97:19]
  wire  ibf_io_in_valid; // @[Frontend.scala 97:19]
  wire [63:0] ibf_io_in_bits_instr; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_in_bits_pc; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[Frontend.scala 97:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[Frontend.scala 97:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[Frontend.scala 97:19]
  wire  ibf_io_out_ready; // @[Frontend.scala 97:19]
  wire  ibf_io_out_valid; // @[Frontend.scala 97:19]
  wire [63:0] ibf_io_out_bits_instr; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_out_bits_pc; // @[Frontend.scala 97:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[Frontend.scala 97:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[Frontend.scala 97:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[Frontend.scala 97:19]
  wire  ibf_io_out_bits_crossPageIPFFix; // @[Frontend.scala 97:19]
  wire  ibf_io_flush; // @[Frontend.scala 97:19]
  wire  idu_clock; // @[Frontend.scala 98:20]
  wire  idu_reset; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_ready; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_valid; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[Frontend.scala 98:20]
  wire  idu_io_in_0_bits_crossPageIPFFix; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_ready; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_valid; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 98:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 98:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 98:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 98:20]
  wire [2:0] idu_io_out_0_bits_ctrl_vtag; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_0_bits_ctrl_vec_addr; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_out_0_bits_ctrl_length_k; // @[Frontend.scala 98:20]
  wire [1:0] idu_io_out_0_bits_ctrl_algorithm; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_ready; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_valid; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_1_bits_cf_instr; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_out_1_bits_cf_pc; // @[Frontend.scala 98:20]
  wire [38:0] idu_io_out_1_bits_cf_pnpc; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_exceptionVec_1; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_exceptionVec_2; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_exceptionVec_12; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_out_1_bits_cf_brIdx; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_cf_crossPageIPFFix; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_ctrl_src1Type; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_ctrl_src2Type; // @[Frontend.scala 98:20]
  wire [2:0] idu_io_out_1_bits_ctrl_fuType; // @[Frontend.scala 98:20]
  wire [6:0] idu_io_out_1_bits_ctrl_fuOpType; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_1_bits_ctrl_rfSrc1; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_1_bits_ctrl_rfSrc2; // @[Frontend.scala 98:20]
  wire  idu_io_out_1_bits_ctrl_rfWen; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_1_bits_ctrl_rfDest; // @[Frontend.scala 98:20]
  wire [2:0] idu_io_out_1_bits_ctrl_vtag; // @[Frontend.scala 98:20]
  wire [4:0] idu_io_out_1_bits_ctrl_vec_addr; // @[Frontend.scala 98:20]
  wire [3:0] idu_io_out_1_bits_ctrl_length_k; // @[Frontend.scala 98:20]
  wire [1:0] idu_io_out_1_bits_ctrl_algorithm; // @[Frontend.scala 98:20]
  wire [63:0] idu_io_out_1_bits_data_imm; // @[Frontend.scala 98:20]
  wire  idu_vmEnable; // @[Frontend.scala 98:20]
  wire [11:0] idu_intrVec; // @[Frontend.scala 98:20]
  wire  FlushableQueue_clock; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_reset; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_enq_valid; // @[FlushableQueue.scala 94:21]
  wire [63:0] FlushableQueue_io_enq_bits_instr; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_enq_bits_pc; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_enq_bits_pnpc; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 94:21]
  wire [3:0] FlushableQueue_io_enq_bits_brIdx; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_deq_ready; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_deq_valid; // @[FlushableQueue.scala 94:21]
  wire [63:0] FlushableQueue_io_deq_bits_instr; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_deq_bits_pc; // @[FlushableQueue.scala 94:21]
  wire [38:0] FlushableQueue_io_deq_bits_pnpc; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_deq_bits_exceptionVec_12; // @[FlushableQueue.scala 94:21]
  wire [3:0] FlushableQueue_io_deq_bits_brIdx; // @[FlushableQueue.scala 94:21]
  wire  FlushableQueue_io_flush; // @[FlushableQueue.scala 94:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [63:0] r_instr; // @[Reg.scala 15:16]
  reg [38:0] r_pc; // @[Reg.scala 15:16]
  reg [38:0] r_pnpc; // @[Reg.scala 15:16]
  reg  r_exceptionVec_12; // @[Reg.scala 15:16]
  reg [3:0] r_brIdx; // @[Reg.scala 15:16]
  reg  r_crossPageIPFFix; // @[Reg.scala 15:16]
  IFU_inorder ifu ( // @[Frontend.scala 96:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ifu_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_ipf(ifu_io_ipf),
    .flushICache(ifu_flushICache),
    .REG_0_valid(ifu_REG_0_valid),
    .REG_0_pc(ifu_REG_0_pc),
    .REG_0_isMissPredict(ifu_REG_0_isMissPredict),
    .REG_0_actualTarget(ifu_REG_0_actualTarget),
    .REG_0_actualTaken(ifu_REG_0_actualTaken),
    .REG_0_fuOpType(ifu_REG_0_fuOpType),
    .REG_0_btbType(ifu_REG_0_btbType),
    .REG_0_isRVC(ifu_REG_0_isRVC),
    .flushTLB(ifu_flushTLB)
  );
  NaiveRVCAlignBuffer ibf ( // @[Frontend.scala 97:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossPageIPFFix(ibf_io_out_bits_crossPageIPFFix),
    .io_flush(ibf_io_flush)
  );
  IDU idu ( // @[Frontend.scala 98:20]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossPageIPFFix(idu_io_in_0_bits_crossPageIPFFix),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(idu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(idu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(idu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(idu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(idu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(idu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(idu_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_cf_runahead_checkpoint_id(idu_io_out_0_bits_cf_runahead_checkpoint_id),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_vtag(idu_io_out_0_bits_ctrl_vtag),
    .io_out_0_bits_ctrl_vec_addr(idu_io_out_0_bits_ctrl_vec_addr),
    .io_out_0_bits_ctrl_length_k(idu_io_out_0_bits_ctrl_length_k),
    .io_out_0_bits_ctrl_algorithm(idu_io_out_0_bits_ctrl_algorithm),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_out_1_ready(idu_io_out_1_ready),
    .io_out_1_valid(idu_io_out_1_valid),
    .io_out_1_bits_cf_instr(idu_io_out_1_bits_cf_instr),
    .io_out_1_bits_cf_pc(idu_io_out_1_bits_cf_pc),
    .io_out_1_bits_cf_pnpc(idu_io_out_1_bits_cf_pnpc),
    .io_out_1_bits_cf_exceptionVec_1(idu_io_out_1_bits_cf_exceptionVec_1),
    .io_out_1_bits_cf_exceptionVec_2(idu_io_out_1_bits_cf_exceptionVec_2),
    .io_out_1_bits_cf_exceptionVec_12(idu_io_out_1_bits_cf_exceptionVec_12),
    .io_out_1_bits_cf_intrVec_0(idu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(idu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(idu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(idu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(idu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(idu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(idu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(idu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(idu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(idu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(idu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(idu_io_out_1_bits_cf_intrVec_11),
    .io_out_1_bits_cf_brIdx(idu_io_out_1_bits_cf_brIdx),
    .io_out_1_bits_cf_crossPageIPFFix(idu_io_out_1_bits_cf_crossPageIPFFix),
    .io_out_1_bits_ctrl_src1Type(idu_io_out_1_bits_ctrl_src1Type),
    .io_out_1_bits_ctrl_src2Type(idu_io_out_1_bits_ctrl_src2Type),
    .io_out_1_bits_ctrl_fuType(idu_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(idu_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_rfSrc1(idu_io_out_1_bits_ctrl_rfSrc1),
    .io_out_1_bits_ctrl_rfSrc2(idu_io_out_1_bits_ctrl_rfSrc2),
    .io_out_1_bits_ctrl_rfWen(idu_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_rfDest(idu_io_out_1_bits_ctrl_rfDest),
    .io_out_1_bits_ctrl_vtag(idu_io_out_1_bits_ctrl_vtag),
    .io_out_1_bits_ctrl_vec_addr(idu_io_out_1_bits_ctrl_vec_addr),
    .io_out_1_bits_ctrl_length_k(idu_io_out_1_bits_ctrl_length_k),
    .io_out_1_bits_ctrl_algorithm(idu_io_out_1_bits_ctrl_algorithm),
    .io_out_1_bits_data_imm(idu_io_out_1_bits_data_imm),
    .vmEnable(idu_vmEnable),
    .intrVec(idu_intrVec)
  );
  FlushableQueue FlushableQueue ( // @[FlushableQueue.scala 94:21]
    .clock(FlushableQueue_clock),
    .reset(FlushableQueue_reset),
    .io_enq_ready(FlushableQueue_io_enq_ready),
    .io_enq_valid(FlushableQueue_io_enq_valid),
    .io_enq_bits_instr(FlushableQueue_io_enq_bits_instr),
    .io_enq_bits_pc(FlushableQueue_io_enq_bits_pc),
    .io_enq_bits_pnpc(FlushableQueue_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_12(FlushableQueue_io_enq_bits_exceptionVec_12),
    .io_enq_bits_brIdx(FlushableQueue_io_enq_bits_brIdx),
    .io_deq_ready(FlushableQueue_io_deq_ready),
    .io_deq_valid(FlushableQueue_io_deq_valid),
    .io_deq_bits_instr(FlushableQueue_io_deq_bits_instr),
    .io_deq_bits_pc(FlushableQueue_io_deq_bits_pc),
    .io_deq_bits_pnpc(FlushableQueue_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_12(FlushableQueue_io_deq_bits_exceptionVec_12),
    .io_deq_bits_brIdx(FlushableQueue_io_deq_bits_brIdx),
    .io_flush(FlushableQueue_io_flush)
  );
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[Frontend.scala 117:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[Frontend.scala 117:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[Frontend.scala 117:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[Frontend.scala 117:11]
  assign io_out_0_valid = idu_io_out_0_valid; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_0 = idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_2 = idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_4 = idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_6 = idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_8 = idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_10 = idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_crossPageIPFFix = idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 112:10]
  assign io_out_0_bits_cf_runahead_checkpoint_id = idu_io_out_0_bits_cf_runahead_checkpoint_id; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_vtag = idu_io_out_0_bits_ctrl_vtag; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_vec_addr = idu_io_out_0_bits_ctrl_vec_addr; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_length_k = idu_io_out_0_bits_ctrl_length_k; // @[Frontend.scala 112:10]
  assign io_out_0_bits_ctrl_algorithm = idu_io_out_0_bits_ctrl_algorithm; // @[Frontend.scala 112:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[Frontend.scala 112:10]
  assign io_out_1_valid = idu_io_out_1_valid; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_instr = idu_io_out_1_bits_cf_instr; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_pc = idu_io_out_1_bits_cf_pc; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_pnpc = idu_io_out_1_bits_cf_pnpc; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_exceptionVec_1 = idu_io_out_1_bits_cf_exceptionVec_1; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_exceptionVec_2 = idu_io_out_1_bits_cf_exceptionVec_2; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_exceptionVec_12 = idu_io_out_1_bits_cf_exceptionVec_12; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_0 = idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_1 = idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_2 = idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_3 = idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_4 = idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_5 = idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_6 = idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_7 = idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_8 = idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_9 = idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_10 = idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_intrVec_11 = idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_brIdx = idu_io_out_1_bits_cf_brIdx; // @[Frontend.scala 112:10]
  assign io_out_1_bits_cf_crossPageIPFFix = idu_io_out_1_bits_cf_crossPageIPFFix; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_src1Type = idu_io_out_1_bits_ctrl_src1Type; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_src2Type = idu_io_out_1_bits_ctrl_src2Type; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_fuType = idu_io_out_1_bits_ctrl_fuType; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_fuOpType = idu_io_out_1_bits_ctrl_fuOpType; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_rfSrc1 = idu_io_out_1_bits_ctrl_rfSrc1; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_rfSrc2 = idu_io_out_1_bits_ctrl_rfSrc2; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_rfWen = idu_io_out_1_bits_ctrl_rfWen; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_rfDest = idu_io_out_1_bits_ctrl_rfDest; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_vtag = idu_io_out_1_bits_ctrl_vtag; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_vec_addr = idu_io_out_1_bits_ctrl_vec_addr; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_length_k = idu_io_out_1_bits_ctrl_length_k; // @[Frontend.scala 112:10]
  assign io_out_1_bits_ctrl_algorithm = idu_io_out_1_bits_ctrl_algorithm; // @[Frontend.scala 112:10]
  assign io_out_1_bits_data_imm = idu_io_out_1_bits_data_imm; // @[Frontend.scala 112:10]
  assign io_flushVec = ifu_io_flushVec; // @[Frontend.scala 114:15]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[Frontend.scala 117:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[Frontend.scala 117:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[Frontend.scala 117:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[Frontend.scala 117:11]
  assign ifu_io_out_ready = FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 98:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[Frontend.scala 113:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[Frontend.scala 113:15]
  assign ifu_io_ipf = io_ipf; // @[Frontend.scala 116:10]
  assign ifu_flushICache = flushICache;
  assign ifu_REG_0_valid = REG_0_valid;
  assign ifu_REG_0_pc = REG_0_pc;
  assign ifu_REG_0_isMissPredict = REG_0_isMissPredict;
  assign ifu_REG_0_actualTarget = REG_0_actualTarget;
  assign ifu_REG_0_actualTaken = REG_0_actualTaken;
  assign ifu_REG_0_fuOpType = REG_0_fuOpType;
  assign ifu_REG_0_btbType = REG_0_btbType;
  assign ifu_REG_0_isRVC = REG_0_isRVC;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = FlushableQueue_io_deq_valid; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_instr = FlushableQueue_io_deq_bits_instr; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_pc = FlushableQueue_io_deq_bits_pc; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_pnpc = FlushableQueue_io_deq_bits_pnpc; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_exceptionVec_12 = FlushableQueue_io_deq_bits_exceptionVec_12; // @[Frontend.scala 104:11]
  assign ibf_io_in_bits_brIdx = FlushableQueue_io_deq_bits_brIdx; // @[Frontend.scala 104:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[Frontend.scala 111:34]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_0_valid = REG; // @[Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = r_instr; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = r_pc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = r_pnpc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = r_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = r_brIdx; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossPageIPFFix = r_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[Frontend.scala 112:10]
  assign idu_io_out_1_ready = io_out_1_ready; // @[Frontend.scala 112:10]
  assign idu_vmEnable = vmEnable;
  assign idu_intrVec = intrVec;
  assign FlushableQueue_clock = clock;
  assign FlushableQueue_reset = reset;
  assign FlushableQueue_io_enq_valid = ifu_io_out_valid; // @[FlushableQueue.scala 95:22]
  assign FlushableQueue_io_enq_bits_instr = ifu_io_out_bits_instr; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_pc = ifu_io_out_bits_pc; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_exceptionVec_12 = ifu_io_out_bits_exceptionVec_12; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[FlushableQueue.scala 96:21]
  assign FlushableQueue_io_deq_ready = ibf_io_in_ready; // @[Frontend.scala 104:11]
  assign FlushableQueue_io_flush = ifu_io_flushVec[0]; // @[Frontend.scala 107:58]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_instr <= ibf_io_out_bits_instr; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_pc <= ibf_io_out_bits_pc; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_pnpc <= ibf_io_out_bits_pnpc; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_brIdx <= ibf_io_out_bits_brIdx; // @[Reg.scala 16:23]
    end
    if (_T_3) begin // @[Reg.scala 16:19]
      r_crossPageIPFFix <= ibf_io_out_bits_crossPageIPFFix; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  r_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  r_exceptionVec_12 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_brIdx = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  r_crossPageIPFFix = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input  [63:0] io_in_0_bits_cf_runahead_checkpoint_id,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input  [2:0]  io_in_0_bits_ctrl_vtag,
  input  [4:0]  io_in_0_bits_ctrl_vec_addr,
  input  [3:0]  io_in_0_bits_ctrl_length_k,
  input  [1:0]  io_in_0_bits_ctrl_algorithm,
  input  [63:0] io_in_0_bits_data_imm,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output [63:0] io_out_bits_cf_runahead_checkpoint_id,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output [2:0]  io_out_bits_ctrl_vtag,
  output [4:0]  io_out_bits_ctrl_vec_addr,
  output [3:0]  io_out_bits_ctrl_length_k,
  output [1:0]  io_out_bits_ctrl_algorithm,
  output [63:0] io_out_bits_data_src1,
  output [63:0] io_out_bits_data_src2,
  output [63:0] io_out_bits_data_imm,
  input         io_wb_rfWen,
  input  [4:0]  io_wb_rfDest,
  input  [63:0] io_wb_rfData,
  input         io_forward_valid,
  input         io_forward_wb_rfWen,
  input  [4:0]  io_forward_wb_rfDest,
  input  [63:0] io_forward_wb_rfData,
  input  [2:0]  io_forward_fuType,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] MEM [0:31]; // @[RF.scala 30:15]
  wire  MEM_MPORT_en; // @[RF.scala 30:15]
  wire [4:0] MEM_MPORT_addr; // @[RF.scala 30:15]
  wire [63:0] MEM_MPORT_data; // @[RF.scala 30:15]
  wire  MEM_MPORT_1_en; // @[RF.scala 30:15]
  wire [4:0] MEM_MPORT_1_addr; // @[RF.scala 30:15]
  wire [63:0] MEM_MPORT_1_data; // @[RF.scala 30:15]
  wire [63:0] MEM_MPORT_2_data; // @[RF.scala 30:15]
  wire [4:0] MEM_MPORT_2_addr; // @[RF.scala 30:15]
  wire  MEM_MPORT_2_mask; // @[RF.scala 30:15]
  wire  MEM_MPORT_2_en; // @[RF.scala 30:15]
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[ISU.scala 43:42]
  wire  dontForward1 = io_forward_fuType != 3'h0 & io_forward_fuType != 3'h1; // @[ISU.scala 44:57]
  wire  src1DependEX = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest &
    forwardRfWen; // @[ISU.scala 41:100]
  wire  src2DependEX = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest &
    forwardRfWen; // @[ISU.scala 41:100]
  wire  src1DependWB = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest & io_wb_rfWen; // @[ISU.scala 41:100]
  wire  src2DependWB = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest & io_wb_rfWen; // @[ISU.scala 41:100]
  wire  _T_14 = ~dontForward1; // @[ISU.scala 50:46]
  wire  src1ForwardNextCycle = src1DependEX & ~dontForward1; // @[ISU.scala 50:43]
  wire  src2ForwardNextCycle = src2DependEX & _T_14; // @[ISU.scala 51:43]
  wire  _T_17 = dontForward1 ? ~src1DependEX : 1'h1; // @[ISU.scala 52:40]
  wire  src1Forward = src1DependWB & _T_17; // @[ISU.scala 52:34]
  wire  _T_19 = dontForward1 ? ~src2DependEX : 1'h1; // @[ISU.scala 53:40]
  wire  src2Forward = src2DependWB & _T_19; // @[ISU.scala 53:34]
  reg [31:0] REG; // @[RF.scala 36:21]
  wire [31:0] _T_20 = REG >> io_in_0_bits_ctrl_rfSrc1; // @[RF.scala 37:37]
  wire  src1Ready = ~_T_20[0] | src1ForwardNextCycle | src1Forward; // @[ISU.scala 56:62]
  wire [31:0] _T_24 = REG >> io_in_0_bits_ctrl_rfSrc2; // @[RF.scala 37:37]
  wire  src2Ready = ~_T_24[0] | src2ForwardNextCycle | src2Forward; // @[ISU.scala 57:62]
  wire [24:0] _T_33 = io_in_0_bits_cf_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_34 = {_T_33,io_in_0_bits_cf_pc}; // @[Cat.scala 30:58]
  wire  _T_35 = ~src1ForwardNextCycle; // @[ISU.scala 66:21]
  wire  _T_36 = src1Forward & ~src1ForwardNextCycle; // @[ISU.scala 66:18]
  wire  _T_41 = ~io_in_0_bits_ctrl_src1Type & _T_35 & ~src1Forward; // @[ISU.scala 67:76]
  wire [63:0] _T_43 = io_in_0_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 : MEM_MPORT_data; // @[RF.scala 31:36]
  wire [63:0] _T_44 = io_in_0_bits_ctrl_src1Type ? _T_34 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_36 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_41 ? _T_43 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_44 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_48 | _T_46; // @[Mux.scala 27:72]
  wire  _T_52 = ~src2ForwardNextCycle; // @[ISU.scala 72:21]
  wire  _T_53 = src2Forward & ~src2ForwardNextCycle; // @[ISU.scala 72:18]
  wire  _T_58 = ~io_in_0_bits_ctrl_src2Type & _T_52 & ~src2Forward; // @[ISU.scala 73:77]
  wire [63:0] _T_60 = io_in_0_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 : MEM_MPORT_1_data; // @[RF.scala 31:36]
  wire [63:0] _T_61 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_62 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_63 = _T_53 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_64 = _T_58 ? _T_60 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_65 = _T_61 | _T_62; // @[Mux.scala 27:72]
  wire [63:0] _T_66 = _T_65 | _T_63; // @[Mux.scala 27:72]
  wire  _T_72 = io_wb_rfDest != 5'h0 & io_wb_rfDest == io_forward_wb_rfDest & forwardRfWen; // @[ISU.scala 41:100]
  wire [62:0] _T_75 = 63'h1 << io_wb_rfDest; // @[RF.scala 38:39]
  wire [31:0] wbClearMask = io_wb_rfWen & ~_T_72 ? _T_75[31:0] : 32'h0; // @[ISU.scala 85:24]
  wire  _T_77 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [62:0] _T_78 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[RF.scala 38:39]
  wire [31:0] isuFireSetMask = _T_77 ? _T_78[31:0] : 32'h0; // @[ISU.scala 87:27]
  wire [31:0] _T_86 = ~wbClearMask; // @[RF.scala 44:26]
  wire [31:0] _T_87 = REG & _T_86; // @[RF.scala 44:24]
  wire [31:0] _T_88 = _T_87 | isuFireSetMask; // @[RF.scala 44:38]
  wire [31:0] _T_90 = {_T_88[31:1],1'h0}; // @[Cat.scala 30:58]
  wire  _T_102 = io_in_0_valid & ~io_out_valid; // @[ISU.scala 101:40]
  wire  _T_105 = io_out_valid & ~_T_77; // @[ISU.scala 102:38]
  wire  _T_106 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign MEM_MPORT_en = 1'h1;
  assign MEM_MPORT_addr = io_in_0_bits_ctrl_rfSrc1;
  assign MEM_MPORT_data = MEM[MEM_MPORT_addr]; // @[RF.scala 30:15]
  assign MEM_MPORT_1_en = 1'h1;
  assign MEM_MPORT_1_addr = io_in_0_bits_ctrl_rfSrc2;
  assign MEM_MPORT_1_data = MEM[MEM_MPORT_1_addr]; // @[RF.scala 30:15]
  assign MEM_MPORT_2_data = io_wb_rfData;
  assign MEM_MPORT_2_addr = io_wb_rfDest;
  assign MEM_MPORT_2_mask = 1'h1;
  assign MEM_MPORT_2_en = io_wb_rfWen;
  assign io_in_0_ready = ~io_in_0_valid | _T_77; // @[ISU.scala 91:37]
  assign io_out_valid = io_in_0_valid & src1Ready & src2Ready; // @[ISU.scala 58:47]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[ISU.scala 77:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[ISU.scala 77:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[ISU.scala 77:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[ISU.scala 77:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[ISU.scala 77:18]
  assign io_out_bits_cf_runahead_checkpoint_id = io_in_0_bits_cf_runahead_checkpoint_id; // @[ISU.scala 77:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[ISU.scala 78:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[ISU.scala 78:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[ISU.scala 78:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[ISU.scala 78:20]
  assign io_out_bits_ctrl_vtag = io_in_0_bits_ctrl_vtag; // @[ISU.scala 78:20]
  assign io_out_bits_ctrl_vec_addr = io_in_0_bits_ctrl_vec_addr; // @[ISU.scala 78:20]
  assign io_out_bits_ctrl_length_k = io_in_0_bits_ctrl_length_k; // @[ISU.scala 78:20]
  assign io_out_bits_ctrl_algorithm = io_in_0_bits_ctrl_algorithm; // @[ISU.scala 78:20]
  assign io_out_bits_data_src1 = _T_49 | _T_47; // @[Mux.scala 27:72]
  assign io_out_bits_data_src2 = _T_66 | _T_64; // @[Mux.scala 27:72]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[ISU.scala 75:25]
  always @(posedge clock) begin
    if (MEM_MPORT_2_en & MEM_MPORT_2_mask) begin
      MEM[MEM_MPORT_2_addr] <= MEM_MPORT_2_data; // @[RF.scala 30:15]
    end
    if (reset) begin // @[RF.scala 36:21]
      REG <= 32'h0; // @[RF.scala 36:21]
    end else if (io_flush) begin // @[ISU.scala 88:19]
      REG <= 32'h0; // @[RF.scala 44:10]
    end else begin
      REG <= _T_90; // @[RF.scala 44:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    MEM[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input  [38:0] io_cfIn_pnpc,
  input  [3:0]  io_cfIn_brIdx,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input  [63:0] io_offset,
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output        REG_0_actualTaken,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[ALU.scala 87:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_in_bits_src2 ^ _T_2; // @[ALU.scala 88:33]
  wire [64:0] _T_4 = io_in_bits_src1 + _T_3; // @[ALU.scala 88:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[ALU.scala 88:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[ALU.scala 88:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[ALU.scala 89:21]
  wire  sltu = ~adderRes[64]; // @[ALU.scala 90:14]
  wire  slt = xorRes[63] ^ sltu; // @[ALU.scala 91:28]
  wire [63:0] _T_10 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_14 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_15 = {_T_14,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_17 = 7'h25 == io_in_bits_func ? _T_10 : io_in_bits_src1; // @[Mux.scala 80:57]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[Mux.scala 80:57]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[ALU.scala 97:18]
  wire [126:0] _GEN_4 = {{63'd0}, shsrc1}; // @[ALU.scala 99:33]
  wire [126:0] _T_23 = _GEN_4 << shamt; // @[ALU.scala 99:33]
  wire [63:0] _T_25 = {63'h0,slt}; // @[Cat.scala 30:58]
  wire [63:0] _T_26 = {63'h0,sltu}; // @[Cat.scala 30:58]
  wire [63:0] _T_27 = shsrc1 >> shamt; // @[ALU.scala 103:32]
  wire [63:0] _T_28 = io_in_bits_src1 | io_in_bits_src2; // @[ALU.scala 104:30]
  wire [63:0] _T_29 = io_in_bits_src1 & io_in_bits_src2; // @[ALU.scala 105:30]
  wire [63:0] _T_30 = 7'h2d == io_in_bits_func ? _T_15 : _T_17; // @[ALU.scala 106:32]
  wire [63:0] _T_32 = $signed(_T_30) >>> shamt; // @[ALU.scala 106:49]
  wire [64:0] _T_34 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _T_23[63:0]} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_36 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _T_25} : _T_34; // @[Mux.scala 80:57]
  wire [64:0] _T_38 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _T_26} : _T_36; // @[Mux.scala 80:57]
  wire [64:0] _T_40 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _T_38; // @[Mux.scala 80:57]
  wire [64:0] _T_42 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _T_27} : _T_40; // @[Mux.scala 80:57]
  wire [64:0] _T_44 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _T_28} : _T_42; // @[Mux.scala 80:57]
  wire [64:0] _T_46 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _T_29} : _T_44; // @[Mux.scala 80:57]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _T_32} : _T_46; // @[Mux.scala 80:57]
  wire [31:0] _T_52 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,res[31:0]}; // @[Cat.scala 30:58]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _T_53} : res; // @[ALU.scala 108:19]
  wire  _T_55 = ~(|xorRes); // @[ALU.scala 111:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[ALU.scala 63:30]
  wire  isBru = io_in_bits_func[4]; // @[ALU.scala 62:31]
  wire  _T_58 = 2'h0 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_59 = 2'h2 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_60 = 2'h3 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_65 = _T_58 & _T_55 | _T_59 & slt | _T_60 & sltu; // @[Mux.scala 27:72]
  wire  taken = _T_65 ^ io_in_bits_func[0]; // @[ALU.scala 118:72]
  wire [63:0] _GEN_1 = {{25'd0}, io_cfIn_pc}; // @[ALU.scala 119:41]
  wire [63:0] _T_68 = _GEN_1 + io_offset; // @[ALU.scala 119:41]
  wire [64:0] _T_69 = isBranch ? {{1'd0}, _T_68} : adderRes; // @[ALU.scala 119:19]
  wire [38:0] target = _T_69[38:0]; // @[ALU.scala 119:63]
  wire  _T_71 = ~taken & isBranch; // @[ALU.scala 120:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[ALU.scala 120:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[ALU.scala 121:35]
  wire [38:0] _T_89 = io_cfIn_pc + 39'h2; // @[ALU.scala 124:71]
  wire [38:0] _T_91 = io_cfIn_pc + 39'h4; // @[ALU.scala 124:89]
  wire [38:0] _T_92 = isRVC ? _T_89 : _T_91; // @[ALU.scala 124:52]
  wire  _T_94 = io_in_valid & isBru; // @[ALU.scala 126:30]
  wire  _T_95 = io_in_valid & isBru & predictWrong; // @[ALU.scala 126:39]
  wire  _T_96 = ~isRVC; // @[ALU.scala 132:33]
  wire [24:0] _T_99 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_100 = {_T_99,io_cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_102 = _T_100 + 64'h4; // @[ALU.scala 132:71]
  wire [63:0] _T_108 = _T_100 + 64'h2; // @[ALU.scala 132:108]
  wire [63:0] _T_109 = ~isRVC ? _T_102 : _T_108; // @[ALU.scala 132:32]
  wire [64:0] _T_110 = isBru ? {{1'd0}, _T_109} : aluRes; // @[ALU.scala 132:21]
  wire  _T_118 = 7'h5c == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_119 = 7'h5e == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_120 = 7'h58 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_121 = 7'h5a == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [1:0] _T_129 = _T_119 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_131 = _T_121 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_2 = {{1'd0}, _T_118}; // @[Mux.scala 27:72]
  wire [1:0] _T_138 = _GEN_2 | _T_129; // @[Mux.scala 27:72]
  wire [1:0] _GEN_3 = {{1'd0}, _T_120}; // @[Mux.scala 27:72]
  wire [1:0] _T_139 = _T_138 | _GEN_3; // @[Mux.scala 27:72]
  reg  REG_valid; // @[ALU.scala 159:34]
  reg [38:0] REG_pc; // @[ALU.scala 159:34]
  reg  REG_isMissPredict; // @[ALU.scala 159:34]
  reg [38:0] REG_actualTarget; // @[ALU.scala 159:34]
  reg  REG_actualTaken; // @[ALU.scala 159:34]
  reg [6:0] REG_fuOpType; // @[ALU.scala 159:34]
  reg [1:0] REG_btbType; // @[ALU.scala 159:34]
  reg  REG_isRVC; // @[ALU.scala 159:34]
  wire  _T_143 = _T_94 & ~predictWrong; // @[ALU.scala 161:32]
  wire  _T_146 = _T_143 & isBranch; // @[ALU.scala 163:33]
  wire  _T_147 = _T_95 & isBranch; // @[ALU.scala 164:33]
  wire  _T_151 = _T_147 & io_cfIn_pc[2:0] == 3'h0; // @[ALU.scala 165:45]
  wire  _T_152 = _T_147 & io_cfIn_pc[2:0] == 3'h0 & isRVC; // @[ALU.scala 165:73]
  wire  _T_158 = _T_151 & _T_96; // @[ALU.scala 166:73]
  wire  _T_162 = _T_147 & io_cfIn_pc[2:0] == 3'h2; // @[ALU.scala 167:45]
  wire  _T_163 = _T_147 & io_cfIn_pc[2:0] == 3'h2 & isRVC; // @[ALU.scala 167:73]
  wire  _T_169 = _T_162 & _T_96; // @[ALU.scala 168:73]
  wire  _T_173 = _T_147 & io_cfIn_pc[2:0] == 3'h4; // @[ALU.scala 169:45]
  wire  _T_174 = _T_147 & io_cfIn_pc[2:0] == 3'h4 & isRVC; // @[ALU.scala 169:73]
  wire  _T_180 = _T_173 & _T_96; // @[ALU.scala 170:73]
  wire  _T_184 = _T_147 & io_cfIn_pc[2:0] == 3'h6; // @[ALU.scala 171:45]
  wire  _T_185 = _T_147 & io_cfIn_pc[2:0] == 3'h6 & isRVC; // @[ALU.scala 171:73]
  wire  _T_191 = _T_184 & _T_96; // @[ALU.scala 172:73]
  wire  _T_194 = io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c; // @[ALU.scala 173:60]
  wire  _T_195 = _T_143 & (io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c); // @[ALU.scala 173:33]
  wire  _T_199 = _T_95 & _T_194; // @[ALU.scala 174:33]
  wire  _T_200 = io_in_bits_func == 7'h5a; // @[ALU.scala 175:41]
  wire  _T_201 = _T_143 & io_in_bits_func == 7'h5a; // @[ALU.scala 175:33]
  wire  _T_203 = _T_95 & _T_200; // @[ALU.scala 176:33]
  wire  _T_204 = io_in_bits_func == 7'h5e; // @[ALU.scala 177:41]
  wire  _T_205 = _T_143 & io_in_bits_func == 7'h5e; // @[ALU.scala 177:33]
  wire  _T_207 = _T_95 & _T_204; // @[ALU.scala 178:33]
  assign io_out_valid = io_in_valid; // @[ALU.scala 146:16]
  assign io_out_bits = _T_110[63:0]; // @[ALU.scala 132:15]
  assign io_redirect_target = _T_71 ? _T_92 : target; // @[ALU.scala 124:28]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[ALU.scala 126:39]
  assign REG_0_valid = REG_valid;
  assign REG_0_pc = REG_pc;
  assign REG_0_isMissPredict = REG_isMissPredict;
  assign REG_0_actualTarget = REG_actualTarget;
  assign REG_0_actualTaken = REG_actualTaken;
  assign REG_0_fuOpType = REG_fuOpType;
  assign REG_0_btbType = REG_btbType;
  assign REG_0_isRVC = REG_isRVC;
  always @(posedge clock) begin
    REG_valid <= io_in_valid & isBru; // @[ALU.scala 149:31]
    REG_pc <= io_cfIn_pc; // @[ALU.scala 159:34]
    if (~taken & isBranch) begin // @[ALU.scala 120:25]
      REG_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      REG_isMissPredict <= ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc;
    end
    REG_actualTarget <= _T_69[38:0]; // @[ALU.scala 119:63]
    REG_actualTaken <= _T_65 ^ io_in_bits_func[0]; // @[ALU.scala 118:72]
    REG_fuOpType <= io_in_bits_func; // @[ALU.scala 159:34]
    REG_btbType <= _T_139 | _T_131; // @[Mux.scala 27:72]
    REG_isRVC <= io_cfIn_instr[1:0] != 2'h3; // @[ALU.scala 121:35]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:122 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[ALU.scala 122:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid | reset)) begin
          $fatal; // @[ALU.scala 122:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG_pc = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  REG_isMissPredict = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  REG_actualTarget = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_actualTaken = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_fuOpType = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  REG_btbType = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  REG_isRVC = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CNNVectorRegFile(
  input         clock,
  input  [4:0]  io_vaddr,
  input  [2:0]  io_vtag,
  input  [2:0]  io_vop,
  input  [3:0]  io_k,
  input         io_vwen,
  input  [79:0] io_load_data,
  input  [39:0] io_load_kernel,
  input  [63:0] io_load_vwidth,
  output [15:0] io_data_main_0,
  output [15:0] io_data_main_1,
  output [15:0] io_data_main_2,
  output [15:0] io_data_main_3,
  output [15:0] io_data_main_4,
  output [15:0] io_data_main_5,
  output [15:0] io_data_main_6,
  output [15:0] io_data_main_7,
  output [15:0] io_data_main_8,
  output [15:0] io_data_main_9,
  output [15:0] io_data_main_10,
  output [15:0] io_data_main_11,
  output [15:0] io_data_main_12,
  output [15:0] io_data_main_13,
  output [15:0] io_data_main_14,
  output [15:0] io_data_main_15,
  output [15:0] io_data_main_16,
  output [15:0] io_data_main_17,
  output [15:0] io_data_main_18,
  output [15:0] io_data_main_19,
  output [15:0] io_data_main_20,
  output [15:0] io_data_main_21,
  output [15:0] io_data_main_22,
  output [15:0] io_data_main_23,
  output [15:0] io_data_main_24,
  output [7:0]  io_data_kernel_0,
  output [7:0]  io_data_kernel_1,
  output [7:0]  io_data_kernel_2,
  output [7:0]  io_data_kernel_3,
  output [7:0]  io_data_kernel_4,
  output [7:0]  io_data_kernel_5,
  output [7:0]  io_data_kernel_6,
  output [7:0]  io_data_kernel_7,
  output [7:0]  io_data_kernel_8,
  output [7:0]  io_data_kernel_9,
  output [7:0]  io_data_kernel_10,
  output [7:0]  io_data_kernel_11,
  output [7:0]  io_data_kernel_12,
  output [7:0]  io_data_kernel_13,
  output [7:0]  io_data_kernel_14,
  output [7:0]  io_data_kernel_15,
  output [7:0]  io_data_kernel_16,
  output [7:0]  io_data_kernel_17,
  output [7:0]  io_data_kernel_18,
  output [7:0]  io_data_kernel_19,
  output [7:0]  io_data_kernel_20,
  output [7:0]  io_data_kernel_21,
  output [7:0]  io_data_kernel_22,
  output [7:0]  io_data_kernel_23,
  output [7:0]  io_data_kernel_24,
  output [3:0]  io_data_kernel_vwidth,
  output [7:0]  io_select_vwidth,
  output [3:0]  io_act_vwidth
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_MEM_INIT
  reg [79:0] vrf_main [0:4]; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_14_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_14_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_14_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_18_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_18_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_18_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_22_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_22_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_22_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_26_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_26_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_26_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_31_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_31_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_31_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_33_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_33_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_33_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_35_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_35_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_35_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_37_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_37_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_37_data; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_39_en; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_39_addr; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_39_data; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_9_data; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_9_addr; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_9_mask; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_9_en; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_13_data; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_13_addr; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_13_mask; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_13_en; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_17_data; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_17_addr; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_17_mask; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_17_en; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_21_data; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_21_addr; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_21_mask; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_21_en; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_25_data; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_25_addr; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_25_mask; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_25_en; // @[CNN_VRF.scala 37:21]
  wire [79:0] vrf_main_MPORT_29_data; // @[CNN_VRF.scala 37:21]
  wire [2:0] vrf_main_MPORT_29_addr; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_29_mask; // @[CNN_VRF.scala 37:21]
  wire  vrf_main_MPORT_29_en; // @[CNN_VRF.scala 37:21]
  reg [39:0] vrf_kernel [0:4]; // @[CNN_VRF.scala 38:23]
  wire  vrf_kernel_MPORT_32_en; // @[CNN_VRF.scala 38:23]
  wire [2:0] vrf_kernel_MPORT_32_addr; // @[CNN_VRF.scala 38:23]
  wire [39:0] vrf_kernel_MPORT_32_data; // @[CNN_VRF.scala 38:23]
  wire  vrf_kernel_MPORT_34_en; // @[CNN_VRF.scala 38:23]
  wire [2:0] vrf_kernel_MPORT_34_addr; // @[CNN_VRF.scala 38:23]
  wire [39:0] vrf_kernel_MPORT_34_data; // @[CNN_VRF.scala 38:23]
  wire  vrf_kernel_MPORT_36_en; // @[CNN_VRF.scala 38:23]
  wire [2:0] vrf_kernel_MPORT_36_addr; // @[CNN_VRF.scala 38:23]
  wire [39:0] vrf_kernel_MPORT_36_data; // @[CNN_VRF.scala 38:23]
  wire  vrf_kernel_MPORT_38_en; // @[CNN_VRF.scala 38:23]
  wire [2:0] vrf_kernel_MPORT_38_addr; // @[CNN_VRF.scala 38:23]
  wire [39:0] vrf_kernel_MPORT_38_data; // @[CNN_VRF.scala 38:23]
  wire  vrf_kernel_MPORT_40_en; // @[CNN_VRF.scala 38:23]
  wire [2:0] vrf_kernel_MPORT_40_addr; // @[CNN_VRF.scala 38:23]
  wire [39:0] vrf_kernel_MPORT_40_data; // @[CNN_VRF.scala 38:23]
  wire [39:0] vrf_kernel_MPORT_11_data; // @[CNN_VRF.scala 38:23]
  wire [2:0] vrf_kernel_MPORT_11_addr; // @[CNN_VRF.scala 38:23]
  wire  vrf_kernel_MPORT_11_mask; // @[CNN_VRF.scala 38:23]
  wire  vrf_kernel_MPORT_11_en; // @[CNN_VRF.scala 38:23]
  reg [3:0] vwidth_kernel [0:4]; // @[CNN_VRF.scala 42:26]
  wire  vwidth_kernel_MPORT_46_en; // @[CNN_VRF.scala 42:26]
  wire [2:0] vwidth_kernel_MPORT_46_addr; // @[CNN_VRF.scala 42:26]
  wire [3:0] vwidth_kernel_MPORT_46_data; // @[CNN_VRF.scala 42:26]
  wire  vwidth_kernel_MPORT_47_en; // @[CNN_VRF.scala 42:26]
  wire [2:0] vwidth_kernel_MPORT_47_addr; // @[CNN_VRF.scala 42:26]
  wire [3:0] vwidth_kernel_MPORT_47_data; // @[CNN_VRF.scala 42:26]
  wire  vwidth_kernel_MPORT_48_en; // @[CNN_VRF.scala 42:26]
  wire [2:0] vwidth_kernel_MPORT_48_addr; // @[CNN_VRF.scala 42:26]
  wire [3:0] vwidth_kernel_MPORT_48_data; // @[CNN_VRF.scala 42:26]
  wire  vwidth_kernel_MPORT_49_en; // @[CNN_VRF.scala 42:26]
  wire [2:0] vwidth_kernel_MPORT_49_addr; // @[CNN_VRF.scala 42:26]
  wire [3:0] vwidth_kernel_MPORT_49_data; // @[CNN_VRF.scala 42:26]
  wire  vwidth_kernel_MPORT_50_en; // @[CNN_VRF.scala 42:26]
  wire [2:0] vwidth_kernel_MPORT_50_addr; // @[CNN_VRF.scala 42:26]
  wire [3:0] vwidth_kernel_MPORT_50_data; // @[CNN_VRF.scala 42:26]
  wire [3:0] vwidth_kernel_MPORT_12_data; // @[CNN_VRF.scala 42:26]
  wire [2:0] vwidth_kernel_MPORT_12_addr; // @[CNN_VRF.scala 42:26]
  wire  vwidth_kernel_MPORT_12_mask; // @[CNN_VRF.scala 42:26]
  wire  vwidth_kernel_MPORT_12_en; // @[CNN_VRF.scala 42:26]
  reg [7:0] global_vwidth [0:7]; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_select_vw_en; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_select_vw_addr; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_select_vw_data; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_en; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_addr; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_data; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_1_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_1_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_1_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_1_en; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_2_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_2_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_2_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_2_en; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_3_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_3_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_3_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_3_en; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_4_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_4_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_4_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_4_en; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_5_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_5_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_5_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_5_en; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_6_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_6_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_6_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_6_en; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_7_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_7_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_7_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_7_en; // @[CNN_VRF.scala 45:26]
  wire [7:0] global_vwidth_MPORT_8_data; // @[CNN_VRF.scala 45:26]
  wire [2:0] global_vwidth_MPORT_8_addr; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_8_mask; // @[CNN_VRF.scala 45:26]
  wire  global_vwidth_MPORT_8_en; // @[CNN_VRF.scala 45:26]
  wire  _T_1 = io_vop == 3'h1; // @[CNN_VRF.scala 49:27]
  wire  vtype = io_vaddr[4]; // @[CNN_VRF.scala 61:23]
  wire  _T_12 = io_vwen & io_vop == 3'h4; // @[CNN_VRF.scala 64:17]
  wire  _T_13 = ~vtype; // @[CNN_VRF.scala 65:19]
  wire  _GEN_26 = ~vtype ? 1'h0 : 1'h1; // @[CNN_VRF.scala 38:23 65:28 69:21]
  wire  _T_18 = io_k >= 4'h1; // @[CNN_VRF.scala 73:18]
  wire  _T_19 = io_k == 4'h1; // @[CNN_VRF.scala 74:35]
  wire  _T_24 = io_k >= 4'h2; // @[CNN_VRF.scala 77:18]
  wire  _T_25 = io_k == 4'h2; // @[CNN_VRF.scala 78:35]
  wire  _T_30 = io_k >= 4'h3; // @[CNN_VRF.scala 81:18]
  wire  _T_31 = io_k == 4'h3; // @[CNN_VRF.scala 82:35]
  wire  _T_36 = io_k >= 4'h4; // @[CNN_VRF.scala 85:18]
  wire  _T_37 = io_k == 4'h4; // @[CNN_VRF.scala 86:35]
  wire  _T_42 = io_k >= 4'h5; // @[CNN_VRF.scala 89:18]
  wire  _GEN_64 = io_vwen & io_vop == 3'h2 & _T_18; // @[CNN_VRF.scala 37:21 72:42]
  wire  _GEN_70 = io_vwen & io_vop == 3'h2 & _T_24; // @[CNN_VRF.scala 37:21 72:42]
  wire  _GEN_76 = io_vwen & io_vop == 3'h2 & _T_30; // @[CNN_VRF.scala 37:21 72:42]
  wire  _GEN_83 = io_vwen & io_vop == 3'h2 & _T_36; // @[CNN_VRF.scala 37:21 72:42]
  wire  _GEN_90 = io_vwen & io_vop == 3'h2 & _T_42; // @[CNN_VRF.scala 37:21 72:42]
  wire [79:0] vrf_main_data_0 = _T_18 ? vrf_main_MPORT_31_data : 80'h0; // @[CNN_VRF.scala 99:32]
  wire [39:0] vrf_kernel_data_0 = _T_18 ? vrf_kernel_MPORT_32_data : 40'h0; // @[CNN_VRF.scala 100:32]
  wire [79:0] vrf_main_data_1 = _T_24 ? vrf_main_MPORT_33_data : 80'h0; // @[CNN_VRF.scala 99:32]
  wire [39:0] vrf_kernel_data_1 = _T_24 ? vrf_kernel_MPORT_34_data : 40'h0; // @[CNN_VRF.scala 100:32]
  wire [79:0] vrf_main_data_2 = _T_30 ? vrf_main_MPORT_35_data : 80'h0; // @[CNN_VRF.scala 99:32]
  wire [39:0] vrf_kernel_data_2 = _T_30 ? vrf_kernel_MPORT_36_data : 40'h0; // @[CNN_VRF.scala 100:32]
  wire [79:0] vrf_main_data_3 = _T_36 ? vrf_main_MPORT_37_data : 80'h0; // @[CNN_VRF.scala 99:32]
  wire [39:0] vrf_kernel_data_3 = _T_36 ? vrf_kernel_MPORT_38_data : 40'h0; // @[CNN_VRF.scala 100:32]
  wire [79:0] vrf_main_data_4 = _T_42 ? vrf_main_MPORT_39_data : 80'h0; // @[CNN_VRF.scala 99:32]
  wire [39:0] vrf_kernel_data_4 = _T_42 ? vrf_kernel_MPORT_40_data : 40'h0; // @[CNN_VRF.scala 100:32]
  wire [3:0] kernel_vw_max_0 = vwidth_kernel_MPORT_46_data; // @[CNN_VRF.scala 116:27 118:35]
  wire [3:0] kernel_vw_max_1 = vwidth_kernel_MPORT_47_data >= kernel_vw_max_0 ? vwidth_kernel_MPORT_47_data :
    kernel_vw_max_0; // @[CNN_VRF.scala 11:8]
  wire [3:0] kernel_vw_max_2 = vwidth_kernel_MPORT_48_data >= kernel_vw_max_1 ? vwidth_kernel_MPORT_48_data :
    kernel_vw_max_1; // @[CNN_VRF.scala 11:8]
  wire [3:0] kernel_vw_max_3 = vwidth_kernel_MPORT_49_data >= kernel_vw_max_2 ? vwidth_kernel_MPORT_49_data :
    kernel_vw_max_2; // @[CNN_VRF.scala 11:8]
  wire [3:0] kernel_vw_max_4 = vwidth_kernel_MPORT_50_data >= kernel_vw_max_3 ? vwidth_kernel_MPORT_50_data :
    kernel_vw_max_3; // @[CNN_VRF.scala 11:8]
  wire [3:0] _T_141 = 4'h1 == io_k ? kernel_vw_max_0 : 4'h0; // @[Mux.scala 80:57]
  wire [3:0] _T_143 = 4'h2 == io_k ? kernel_vw_max_1 : _T_141; // @[Mux.scala 80:57]
  wire [3:0] _T_145 = 4'h3 == io_k ? kernel_vw_max_2 : _T_143; // @[Mux.scala 80:57]
  wire [3:0] _T_147 = 4'h4 == io_k ? kernel_vw_max_3 : _T_145; // @[Mux.scala 80:57]
  assign vrf_main_MPORT_14_en = _T_12 ? 1'h0 : _GEN_64;
  assign vrf_main_MPORT_14_addr = 3'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_14_data = vrf_main[vrf_main_MPORT_14_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_14_data = vrf_main_MPORT_14_addr >= 3'h5 ? _RAND_1[79:0] : vrf_main[vrf_main_MPORT_14_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_18_en = _T_12 ? 1'h0 : _GEN_70;
  assign vrf_main_MPORT_18_addr = 3'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_18_data = vrf_main[vrf_main_MPORT_18_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_18_data = vrf_main_MPORT_18_addr >= 3'h5 ? _RAND_2[79:0] : vrf_main[vrf_main_MPORT_18_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_22_en = _T_12 ? 1'h0 : _GEN_76;
  assign vrf_main_MPORT_22_addr = 3'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_22_data = vrf_main[vrf_main_MPORT_22_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_22_data = vrf_main_MPORT_22_addr >= 3'h5 ? _RAND_3[79:0] : vrf_main[vrf_main_MPORT_22_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_26_en = _T_12 ? 1'h0 : _GEN_83;
  assign vrf_main_MPORT_26_addr = 3'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_26_data = vrf_main[vrf_main_MPORT_26_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_26_data = vrf_main_MPORT_26_addr >= 3'h5 ? _RAND_4[79:0] : vrf_main[vrf_main_MPORT_26_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_31_en = 1'h1;
  assign vrf_main_MPORT_31_addr = 3'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_31_data = vrf_main[vrf_main_MPORT_31_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_31_data = vrf_main_MPORT_31_addr >= 3'h5 ? _RAND_5[79:0] : vrf_main[vrf_main_MPORT_31_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_33_en = 1'h1;
  assign vrf_main_MPORT_33_addr = 3'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_33_data = vrf_main[vrf_main_MPORT_33_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_33_data = vrf_main_MPORT_33_addr >= 3'h5 ? _RAND_6[79:0] : vrf_main[vrf_main_MPORT_33_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_35_en = 1'h1;
  assign vrf_main_MPORT_35_addr = 3'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_35_data = vrf_main[vrf_main_MPORT_35_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_35_data = vrf_main_MPORT_35_addr >= 3'h5 ? _RAND_7[79:0] : vrf_main[vrf_main_MPORT_35_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_37_en = 1'h1;
  assign vrf_main_MPORT_37_addr = 3'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_37_data = vrf_main[vrf_main_MPORT_37_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_37_data = vrf_main_MPORT_37_addr >= 3'h5 ? _RAND_8[79:0] : vrf_main[vrf_main_MPORT_37_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_39_en = 1'h1;
  assign vrf_main_MPORT_39_addr = 3'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_39_data = vrf_main[vrf_main_MPORT_39_addr]; // @[CNN_VRF.scala 37:21]
  `else
  assign vrf_main_MPORT_39_data = vrf_main_MPORT_39_addr >= 3'h5 ? _RAND_9[79:0] : vrf_main[vrf_main_MPORT_39_addr]; // @[CNN_VRF.scala 37:21]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_main_MPORT_9_data = io_load_data;
  assign vrf_main_MPORT_9_addr = io_vaddr[2:0];
  assign vrf_main_MPORT_9_mask = 1'h1;
  assign vrf_main_MPORT_9_en = _T_12 & _T_13;
  assign vrf_main_MPORT_13_data = _T_19 ? io_load_data : vrf_main_MPORT_14_data;
  assign vrf_main_MPORT_13_addr = 3'h0;
  assign vrf_main_MPORT_13_mask = 1'h1;
  assign vrf_main_MPORT_13_en = _T_12 ? 1'h0 : _GEN_64;
  assign vrf_main_MPORT_17_data = _T_25 ? io_load_data : vrf_main_MPORT_18_data;
  assign vrf_main_MPORT_17_addr = 3'h1;
  assign vrf_main_MPORT_17_mask = 1'h1;
  assign vrf_main_MPORT_17_en = _T_12 ? 1'h0 : _GEN_70;
  assign vrf_main_MPORT_21_data = _T_31 ? io_load_data : vrf_main_MPORT_22_data;
  assign vrf_main_MPORT_21_addr = 3'h2;
  assign vrf_main_MPORT_21_mask = 1'h1;
  assign vrf_main_MPORT_21_en = _T_12 ? 1'h0 : _GEN_76;
  assign vrf_main_MPORT_25_data = _T_37 ? io_load_data : vrf_main_MPORT_26_data;
  assign vrf_main_MPORT_25_addr = 3'h3;
  assign vrf_main_MPORT_25_mask = 1'h1;
  assign vrf_main_MPORT_25_en = _T_12 ? 1'h0 : _GEN_83;
  assign vrf_main_MPORT_29_data = io_load_data;
  assign vrf_main_MPORT_29_addr = 3'h4;
  assign vrf_main_MPORT_29_mask = 1'h1;
  assign vrf_main_MPORT_29_en = _T_12 ? 1'h0 : _GEN_90;
  assign vrf_kernel_MPORT_32_en = 1'h1;
  assign vrf_kernel_MPORT_32_addr = 3'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_32_data = vrf_kernel[vrf_kernel_MPORT_32_addr]; // @[CNN_VRF.scala 38:23]
  `else
  assign vrf_kernel_MPORT_32_data = vrf_kernel_MPORT_32_addr >= 3'h5 ? _RAND_11[39:0] :
    vrf_kernel[vrf_kernel_MPORT_32_addr]; // @[CNN_VRF.scala 38:23]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_34_en = 1'h1;
  assign vrf_kernel_MPORT_34_addr = 3'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_34_data = vrf_kernel[vrf_kernel_MPORT_34_addr]; // @[CNN_VRF.scala 38:23]
  `else
  assign vrf_kernel_MPORT_34_data = vrf_kernel_MPORT_34_addr >= 3'h5 ? _RAND_12[39:0] :
    vrf_kernel[vrf_kernel_MPORT_34_addr]; // @[CNN_VRF.scala 38:23]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_36_en = 1'h1;
  assign vrf_kernel_MPORT_36_addr = 3'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_36_data = vrf_kernel[vrf_kernel_MPORT_36_addr]; // @[CNN_VRF.scala 38:23]
  `else
  assign vrf_kernel_MPORT_36_data = vrf_kernel_MPORT_36_addr >= 3'h5 ? _RAND_13[39:0] :
    vrf_kernel[vrf_kernel_MPORT_36_addr]; // @[CNN_VRF.scala 38:23]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_38_en = 1'h1;
  assign vrf_kernel_MPORT_38_addr = 3'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_38_data = vrf_kernel[vrf_kernel_MPORT_38_addr]; // @[CNN_VRF.scala 38:23]
  `else
  assign vrf_kernel_MPORT_38_data = vrf_kernel_MPORT_38_addr >= 3'h5 ? _RAND_14[39:0] :
    vrf_kernel[vrf_kernel_MPORT_38_addr]; // @[CNN_VRF.scala 38:23]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_40_en = 1'h1;
  assign vrf_kernel_MPORT_40_addr = 3'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_40_data = vrf_kernel[vrf_kernel_MPORT_40_addr]; // @[CNN_VRF.scala 38:23]
  `else
  assign vrf_kernel_MPORT_40_data = vrf_kernel_MPORT_40_addr >= 3'h5 ? _RAND_15[39:0] :
    vrf_kernel[vrf_kernel_MPORT_40_addr]; // @[CNN_VRF.scala 38:23]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vrf_kernel_MPORT_11_data = io_load_kernel;
  assign vrf_kernel_MPORT_11_addr = io_vaddr[2:0];
  assign vrf_kernel_MPORT_11_mask = 1'h1;
  assign vrf_kernel_MPORT_11_en = _T_12 & _GEN_26;
  assign vwidth_kernel_MPORT_46_en = 1'h1;
  assign vwidth_kernel_MPORT_46_addr = 3'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_46_data = vwidth_kernel[vwidth_kernel_MPORT_46_addr]; // @[CNN_VRF.scala 42:26]
  `else
  assign vwidth_kernel_MPORT_46_data = vwidth_kernel_MPORT_46_addr >= 3'h5 ? _RAND_17[3:0] :
    vwidth_kernel[vwidth_kernel_MPORT_46_addr]; // @[CNN_VRF.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_47_en = 1'h1;
  assign vwidth_kernel_MPORT_47_addr = 3'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_47_data = vwidth_kernel[vwidth_kernel_MPORT_47_addr]; // @[CNN_VRF.scala 42:26]
  `else
  assign vwidth_kernel_MPORT_47_data = vwidth_kernel_MPORT_47_addr >= 3'h5 ? _RAND_18[3:0] :
    vwidth_kernel[vwidth_kernel_MPORT_47_addr]; // @[CNN_VRF.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_48_en = 1'h1;
  assign vwidth_kernel_MPORT_48_addr = 3'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_48_data = vwidth_kernel[vwidth_kernel_MPORT_48_addr]; // @[CNN_VRF.scala 42:26]
  `else
  assign vwidth_kernel_MPORT_48_data = vwidth_kernel_MPORT_48_addr >= 3'h5 ? _RAND_19[3:0] :
    vwidth_kernel[vwidth_kernel_MPORT_48_addr]; // @[CNN_VRF.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_49_en = 1'h1;
  assign vwidth_kernel_MPORT_49_addr = 3'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_49_data = vwidth_kernel[vwidth_kernel_MPORT_49_addr]; // @[CNN_VRF.scala 42:26]
  `else
  assign vwidth_kernel_MPORT_49_data = vwidth_kernel_MPORT_49_addr >= 3'h5 ? _RAND_20[3:0] :
    vwidth_kernel[vwidth_kernel_MPORT_49_addr]; // @[CNN_VRF.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_50_en = 1'h1;
  assign vwidth_kernel_MPORT_50_addr = 3'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_50_data = vwidth_kernel[vwidth_kernel_MPORT_50_addr]; // @[CNN_VRF.scala 42:26]
  `else
  assign vwidth_kernel_MPORT_50_data = vwidth_kernel_MPORT_50_addr >= 3'h5 ? _RAND_21[3:0] :
    vwidth_kernel[vwidth_kernel_MPORT_50_addr]; // @[CNN_VRF.scala 42:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign vwidth_kernel_MPORT_12_data = global_vwidth_select_vw_data[3:0];
  assign vwidth_kernel_MPORT_12_addr = io_vaddr[2:0];
  assign vwidth_kernel_MPORT_12_mask = 1'h1;
  assign vwidth_kernel_MPORT_12_en = _T_12 & _GEN_26;
  assign global_vwidth_select_vw_en = 1'h1;
  assign global_vwidth_select_vw_addr = io_vtag;
  assign global_vwidth_select_vw_data = global_vwidth[global_vwidth_select_vw_addr]; // @[CNN_VRF.scala 45:26]
  assign global_vwidth_MPORT_en = 1'h1;
  assign global_vwidth_MPORT_addr = 3'h0;
  assign global_vwidth_MPORT_data = global_vwidth[global_vwidth_MPORT_addr]; // @[CNN_VRF.scala 45:26]
  assign global_vwidth_MPORT_1_data = io_load_vwidth[7:0];
  assign global_vwidth_MPORT_1_addr = 3'h0;
  assign global_vwidth_MPORT_1_mask = 1'h1;
  assign global_vwidth_MPORT_1_en = io_vwen & _T_1;
  assign global_vwidth_MPORT_2_data = io_load_vwidth[15:8];
  assign global_vwidth_MPORT_2_addr = 3'h1;
  assign global_vwidth_MPORT_2_mask = 1'h1;
  assign global_vwidth_MPORT_2_en = io_vwen & _T_1;
  assign global_vwidth_MPORT_3_data = io_load_vwidth[23:16];
  assign global_vwidth_MPORT_3_addr = 3'h2;
  assign global_vwidth_MPORT_3_mask = 1'h1;
  assign global_vwidth_MPORT_3_en = io_vwen & _T_1;
  assign global_vwidth_MPORT_4_data = io_load_vwidth[31:24];
  assign global_vwidth_MPORT_4_addr = 3'h3;
  assign global_vwidth_MPORT_4_mask = 1'h1;
  assign global_vwidth_MPORT_4_en = io_vwen & _T_1;
  assign global_vwidth_MPORT_5_data = io_load_vwidth[39:32];
  assign global_vwidth_MPORT_5_addr = 3'h4;
  assign global_vwidth_MPORT_5_mask = 1'h1;
  assign global_vwidth_MPORT_5_en = io_vwen & _T_1;
  assign global_vwidth_MPORT_6_data = io_load_vwidth[47:40];
  assign global_vwidth_MPORT_6_addr = 3'h5;
  assign global_vwidth_MPORT_6_mask = 1'h1;
  assign global_vwidth_MPORT_6_en = io_vwen & _T_1;
  assign global_vwidth_MPORT_7_data = io_load_vwidth[55:48];
  assign global_vwidth_MPORT_7_addr = 3'h6;
  assign global_vwidth_MPORT_7_mask = 1'h1;
  assign global_vwidth_MPORT_7_en = io_vwen & _T_1;
  assign global_vwidth_MPORT_8_data = io_load_vwidth[63:56];
  assign global_vwidth_MPORT_8_addr = 3'h7;
  assign global_vwidth_MPORT_8_mask = 1'h1;
  assign global_vwidth_MPORT_8_en = io_vwen & _T_1;
  assign io_data_main_0 = vrf_main_data_0[15:0]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_1 = vrf_main_data_1[15:0]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_2 = vrf_main_data_2[15:0]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_3 = vrf_main_data_3[15:0]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_4 = vrf_main_data_4[15:0]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_5 = vrf_main_data_0[31:16]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_6 = vrf_main_data_1[31:16]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_7 = vrf_main_data_2[31:16]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_8 = vrf_main_data_3[31:16]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_9 = vrf_main_data_4[31:16]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_10 = vrf_main_data_0[47:32]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_11 = vrf_main_data_1[47:32]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_12 = vrf_main_data_2[47:32]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_13 = vrf_main_data_3[47:32]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_14 = vrf_main_data_4[47:32]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_15 = vrf_main_data_0[63:48]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_16 = vrf_main_data_1[63:48]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_17 = vrf_main_data_2[63:48]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_18 = vrf_main_data_3[63:48]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_19 = vrf_main_data_4[63:48]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_20 = vrf_main_data_0[79:64]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_21 = vrf_main_data_1[79:64]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_22 = vrf_main_data_2[79:64]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_23 = vrf_main_data_3[79:64]; // @[CNN_VRF.scala 105:52]
  assign io_data_main_24 = vrf_main_data_4[79:64]; // @[CNN_VRF.scala 105:52]
  assign io_data_kernel_0 = vrf_kernel_data_0[7:0]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_1 = vrf_kernel_data_0[15:8]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_2 = vrf_kernel_data_0[23:16]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_3 = vrf_kernel_data_0[31:24]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_4 = vrf_kernel_data_0[39:32]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_5 = vrf_kernel_data_1[7:0]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_6 = vrf_kernel_data_1[15:8]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_7 = vrf_kernel_data_1[23:16]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_8 = vrf_kernel_data_1[31:24]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_9 = vrf_kernel_data_1[39:32]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_10 = vrf_kernel_data_2[7:0]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_11 = vrf_kernel_data_2[15:8]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_12 = vrf_kernel_data_2[23:16]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_13 = vrf_kernel_data_2[31:24]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_14 = vrf_kernel_data_2[39:32]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_15 = vrf_kernel_data_3[7:0]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_16 = vrf_kernel_data_3[15:8]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_17 = vrf_kernel_data_3[23:16]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_18 = vrf_kernel_data_3[31:24]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_19 = vrf_kernel_data_3[39:32]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_20 = vrf_kernel_data_4[7:0]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_21 = vrf_kernel_data_4[15:8]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_22 = vrf_kernel_data_4[23:16]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_23 = vrf_kernel_data_4[31:24]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_24 = vrf_kernel_data_4[39:32]; // @[CNN_VRF.scala 106:54]
  assign io_data_kernel_vwidth = 4'h5 == io_k ? kernel_vw_max_4 : _T_147; // @[Mux.scala 80:57]
  assign io_select_vwidth = global_vwidth_select_vw_data; // @[CNN_VRF.scala 47:20]
  assign io_act_vwidth = global_vwidth_MPORT_data[7:4]; // @[CNN_VRF.scala 48:36]
  always @(posedge clock) begin
    if (vrf_main_MPORT_9_en & vrf_main_MPORT_9_mask) begin
      vrf_main[vrf_main_MPORT_9_addr] <= vrf_main_MPORT_9_data; // @[CNN_VRF.scala 37:21]
    end
    if (vrf_main_MPORT_13_en & vrf_main_MPORT_13_mask) begin
      vrf_main[vrf_main_MPORT_13_addr] <= vrf_main_MPORT_13_data; // @[CNN_VRF.scala 37:21]
    end
    if (vrf_main_MPORT_17_en & vrf_main_MPORT_17_mask) begin
      vrf_main[vrf_main_MPORT_17_addr] <= vrf_main_MPORT_17_data; // @[CNN_VRF.scala 37:21]
    end
    if (vrf_main_MPORT_21_en & vrf_main_MPORT_21_mask) begin
      vrf_main[vrf_main_MPORT_21_addr] <= vrf_main_MPORT_21_data; // @[CNN_VRF.scala 37:21]
    end
    if (vrf_main_MPORT_25_en & vrf_main_MPORT_25_mask) begin
      vrf_main[vrf_main_MPORT_25_addr] <= vrf_main_MPORT_25_data; // @[CNN_VRF.scala 37:21]
    end
    if (vrf_main_MPORT_29_en & vrf_main_MPORT_29_mask) begin
      vrf_main[vrf_main_MPORT_29_addr] <= vrf_main_MPORT_29_data; // @[CNN_VRF.scala 37:21]
    end
    if (vrf_kernel_MPORT_11_en & vrf_kernel_MPORT_11_mask) begin
      vrf_kernel[vrf_kernel_MPORT_11_addr] <= vrf_kernel_MPORT_11_data; // @[CNN_VRF.scala 38:23]
    end
    if (vwidth_kernel_MPORT_12_en & vwidth_kernel_MPORT_12_mask) begin
      vwidth_kernel[vwidth_kernel_MPORT_12_addr] <= vwidth_kernel_MPORT_12_data; // @[CNN_VRF.scala 42:26]
    end
    if (global_vwidth_MPORT_1_en & global_vwidth_MPORT_1_mask) begin
      global_vwidth[global_vwidth_MPORT_1_addr] <= global_vwidth_MPORT_1_data; // @[CNN_VRF.scala 45:26]
    end
    if (global_vwidth_MPORT_2_en & global_vwidth_MPORT_2_mask) begin
      global_vwidth[global_vwidth_MPORT_2_addr] <= global_vwidth_MPORT_2_data; // @[CNN_VRF.scala 45:26]
    end
    if (global_vwidth_MPORT_3_en & global_vwidth_MPORT_3_mask) begin
      global_vwidth[global_vwidth_MPORT_3_addr] <= global_vwidth_MPORT_3_data; // @[CNN_VRF.scala 45:26]
    end
    if (global_vwidth_MPORT_4_en & global_vwidth_MPORT_4_mask) begin
      global_vwidth[global_vwidth_MPORT_4_addr] <= global_vwidth_MPORT_4_data; // @[CNN_VRF.scala 45:26]
    end
    if (global_vwidth_MPORT_5_en & global_vwidth_MPORT_5_mask) begin
      global_vwidth[global_vwidth_MPORT_5_addr] <= global_vwidth_MPORT_5_data; // @[CNN_VRF.scala 45:26]
    end
    if (global_vwidth_MPORT_6_en & global_vwidth_MPORT_6_mask) begin
      global_vwidth[global_vwidth_MPORT_6_addr] <= global_vwidth_MPORT_6_data; // @[CNN_VRF.scala 45:26]
    end
    if (global_vwidth_MPORT_7_en & global_vwidth_MPORT_7_mask) begin
      global_vwidth[global_vwidth_MPORT_7_addr] <= global_vwidth_MPORT_7_data; // @[CNN_VRF.scala 45:26]
    end
    if (global_vwidth_MPORT_8_en & global_vwidth_MPORT_8_mask) begin
      global_vwidth[global_vwidth_MPORT_8_addr] <= global_vwidth_MPORT_8_data; // @[CNN_VRF.scala 45:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {3{`RANDOM}};
  _RAND_2 = {3{`RANDOM}};
  _RAND_3 = {3{`RANDOM}};
  _RAND_4 = {3{`RANDOM}};
  _RAND_5 = {3{`RANDOM}};
  _RAND_6 = {3{`RANDOM}};
  _RAND_7 = {3{`RANDOM}};
  _RAND_8 = {3{`RANDOM}};
  _RAND_9 = {3{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
  _RAND_12 = {2{`RANDOM}};
  _RAND_13 = {2{`RANDOM}};
  _RAND_14 = {2{`RANDOM}};
  _RAND_15 = {2{`RANDOM}};
  _RAND_17 = {1{`RANDOM}};
  _RAND_18 = {1{`RANDOM}};
  _RAND_19 = {1{`RANDOM}};
  _RAND_20 = {1{`RANDOM}};
  _RAND_21 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    vrf_main[initvar] = _RAND_0[79:0];
  _RAND_10 = {2{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    vrf_kernel[initvar] = _RAND_10[39:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    vwidth_kernel[initvar] = _RAND_16[3:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    global_vwidth[initvar] = _RAND_22[7:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoothEncoderP(
  input  [2:0]  io_y,
  input  [31:0] io_x,
  output [31:0] io_p
);
  wire [32:0] _T = {io_x, 1'h0}; // @[CNN_CONV.scala 21:23]
  wire [32:0] _T_2 = ~_T; // @[CNN_CONV.scala 22:17]
  wire [31:0] _T_3 = ~io_x; // @[CNN_CONV.scala 23:17]
  wire  _T_6 = 3'h1 == io_y; // @[LookupTree.scala 24:34]
  wire  _T_7 = 3'h2 == io_y; // @[LookupTree.scala 24:34]
  wire  _T_8 = 3'h3 == io_y; // @[LookupTree.scala 24:34]
  wire  _T_9 = 3'h4 == io_y; // @[LookupTree.scala 24:34]
  wire  _T_10 = 3'h5 == io_y; // @[LookupTree.scala 24:34]
  wire  _T_11 = 3'h6 == io_y; // @[LookupTree.scala 24:34]
  wire [31:0] _T_14 = _T_6 ? io_x : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_15 = _T_7 ? io_x : 32'h0; // @[Mux.scala 27:72]
  wire [32:0] _T_16 = _T_8 ? _T : 33'h0; // @[Mux.scala 27:72]
  wire [32:0] _T_17 = _T_9 ? _T_2 : 33'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_18 = _T_10 ? _T_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_19 = _T_11 ? _T_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_22 = _T_14 | _T_15; // @[Mux.scala 27:72]
  wire [32:0] _GEN_0 = {{1'd0}, _T_22}; // @[Mux.scala 27:72]
  wire [32:0] _T_23 = _GEN_0 | _T_16; // @[Mux.scala 27:72]
  wire [32:0] _T_24 = _T_23 | _T_17; // @[Mux.scala 27:72]
  wire [32:0] _GEN_1 = {{1'd0}, _T_18}; // @[Mux.scala 27:72]
  wire [32:0] _T_25 = _T_24 | _GEN_1; // @[Mux.scala 27:72]
  wire [32:0] _GEN_2 = {{1'd0}, _T_19}; // @[Mux.scala 27:72]
  wire [32:0] _T_26 = _T_25 | _GEN_2; // @[Mux.scala 27:72]
  assign io_p = _T_26[31:0]; // @[CNN_CONV.scala 17:8]
endmodule
module BoothEncoderC(
  input  [2:0] io_y,
  output       io_c
);
  assign io_c = 3'h6 == io_y | (3'h5 == io_y | 3'h4 == io_y); // @[Mux.scala 80:57]
endmodule
module WallaceTree25(
  input  [24:0] io_n,
  input  [23:0] io_cin,
  output        io_s,
  output        io_c,
  output [23:0] io_cout
);
  wire  ly1_out_0 = io_n[0] ^ io_n[1] ^ io_n[2]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_0 = io_n[0] & io_n[1] | io_n[0] & io_n[2] | io_n[1] & io_n[2]; // @[CNN_CONV.scala 64:21]
  wire  ly1_out_1 = io_n[3] ^ io_n[4] ^ io_n[5]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_1 = io_n[3] & io_n[4] | io_n[3] & io_n[5] | io_n[4] & io_n[5]; // @[CNN_CONV.scala 64:21]
  wire  ly1_out_2 = io_n[6] ^ io_n[7] ^ io_n[8]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_2 = io_n[6] & io_n[7] | io_n[6] & io_n[8] | io_n[7] & io_n[8]; // @[CNN_CONV.scala 64:21]
  wire  ly1_out_3 = io_n[9] ^ io_n[10] ^ io_n[11]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_3 = io_n[9] & io_n[10] | io_n[9] & io_n[11] | io_n[10] & io_n[11]; // @[CNN_CONV.scala 64:21]
  wire  ly1_out_4 = io_n[12] ^ io_n[13] ^ io_n[14]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_4 = io_n[12] & io_n[13] | io_n[12] & io_n[14] | io_n[13] & io_n[14]; // @[CNN_CONV.scala 64:21]
  wire  ly1_out_5 = io_n[15] ^ io_n[16] ^ io_n[17]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_5 = io_n[15] & io_n[16] | io_n[15] & io_n[17] | io_n[16] & io_n[17]; // @[CNN_CONV.scala 64:21]
  wire  ly1_out_6 = io_n[18] ^ io_n[19] ^ io_n[20]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_6 = io_n[18] & io_n[19] | io_n[18] & io_n[20] | io_n[19] & io_n[20]; // @[CNN_CONV.scala 64:21]
  wire  ly1_out_7 = io_n[21] ^ io_n[22] ^ io_n[23]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_7 = io_n[21] & io_n[22] | io_n[21] & io_n[23] | io_n[22] & io_n[23]; // @[CNN_CONV.scala 64:21]
  wire [16:0] ly2_in = {ly1_out_7,ly1_out_6,ly1_out_5,ly1_out_4,ly1_out_3,ly1_out_2,ly1_out_1,ly1_out_0,io_cin[7:0],io_n
    [24]}; // @[Cat.scala 30:58]
  wire  ly2_out_0 = ly2_in[0] ^ ly2_in[1] ^ ly2_in[2]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_8 = ly2_in[0] & ly2_in[1] | ly2_in[0] & ly2_in[2] | ly2_in[1] & ly2_in[2]; // @[CNN_CONV.scala 64:21]
  wire  ly2_out_1 = ly2_in[3] ^ ly2_in[4] ^ ly2_in[5]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_9 = ly2_in[3] & ly2_in[4] | ly2_in[3] & ly2_in[5] | ly2_in[4] & ly2_in[5]; // @[CNN_CONV.scala 64:21]
  wire  ly2_out_2 = ly2_in[6] ^ ly2_in[7] ^ ly2_in[8]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_10 = ly2_in[6] & ly2_in[7] | ly2_in[6] & ly2_in[8] | ly2_in[7] & ly2_in[8]; // @[CNN_CONV.scala 64:21]
  wire  ly2_out_3 = ly2_in[9] ^ ly2_in[10] ^ ly2_in[11]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_11 = ly2_in[9] & ly2_in[10] | ly2_in[9] & ly2_in[11] | ly2_in[10] & ly2_in[11]; // @[CNN_CONV.scala 64:21]
  wire  ly2_out_4 = ly2_in[12] ^ ly2_in[13] ^ ly2_in[14]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_12 = ly2_in[12] & ly2_in[13] | ly2_in[12] & ly2_in[14] | ly2_in[13] & ly2_in[14]; // @[CNN_CONV.scala 64:21]
  wire  ly2_out_5 = ly2_in[15] ^ ly2_in[16]; // @[CNN_CONV.scala 69:7]
  wire  out_cout_13 = ly2_in[15] & ly2_in[16]; // @[CNN_CONV.scala 74:7]
  wire [11:0] ly3_in = {ly2_out_5,ly2_out_4,ly2_out_3,ly2_out_2,ly2_out_1,ly2_out_0,io_cin[13:8]}; // @[Cat.scala 30:58]
  wire  ly3_out_0 = ly3_in[0] ^ ly3_in[1] ^ ly3_in[2]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_14 = ly3_in[0] & ly3_in[1] | ly3_in[0] & ly3_in[2] | ly3_in[1] & ly3_in[2]; // @[CNN_CONV.scala 64:21]
  wire  ly3_out_1 = ly3_in[3] ^ ly3_in[4] ^ ly3_in[5]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_15 = ly3_in[3] & ly3_in[4] | ly3_in[3] & ly3_in[5] | ly3_in[4] & ly3_in[5]; // @[CNN_CONV.scala 64:21]
  wire  ly3_out_2 = ly3_in[6] ^ ly3_in[7] ^ ly3_in[8]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_16 = ly3_in[6] & ly3_in[7] | ly3_in[6] & ly3_in[8] | ly3_in[7] & ly3_in[8]; // @[CNN_CONV.scala 64:21]
  wire  ly3_out_3 = ly3_in[9] ^ ly3_in[10] ^ ly3_in[11]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_17 = ly3_in[9] & ly3_in[10] | ly3_in[9] & ly3_in[11] | ly3_in[10] & ly3_in[11]; // @[CNN_CONV.scala 64:21]
  wire [7:0] ly4_in = {ly3_out_3,ly3_out_2,ly3_out_1,ly3_out_0,io_cin[17:14]}; // @[Cat.scala 30:58]
  wire  ly4_out_0 = ly4_in[0] ^ ly4_in[1] ^ ly4_in[2]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_18 = ly4_in[0] & ly4_in[1] | ly4_in[0] & ly4_in[2] | ly4_in[1] & ly4_in[2]; // @[CNN_CONV.scala 64:21]
  wire  ly4_out_1 = ly4_in[3] ^ ly4_in[4] ^ ly4_in[5]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_19 = ly4_in[3] & ly4_in[4] | ly4_in[3] & ly4_in[5] | ly4_in[4] & ly4_in[5]; // @[CNN_CONV.scala 64:21]
  wire  ly4_out_2 = ly4_in[6] ^ ly4_in[7]; // @[CNN_CONV.scala 69:7]
  wire  out_cout_20 = ly4_in[6] & ly4_in[7]; // @[CNN_CONV.scala 74:7]
  wire [5:0] ly5_in = {ly4_out_2,ly4_out_1,ly4_out_0,io_cin[20:18]}; // @[Cat.scala 30:58]
  wire  ly5_out_0 = ly5_in[0] ^ ly5_in[1] ^ ly5_in[2]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_21 = ly5_in[0] & ly5_in[1] | ly5_in[0] & ly5_in[2] | ly5_in[1] & ly5_in[2]; // @[CNN_CONV.scala 64:21]
  wire  ly5_out_1 = ly5_in[3] ^ ly5_in[4] ^ ly5_in[5]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_22 = ly5_in[3] & ly5_in[4] | ly5_in[3] & ly5_in[5] | ly5_in[4] & ly5_in[5]; // @[CNN_CONV.scala 64:21]
  wire [2:0] ly6_in = {ly5_out_1,ly5_out_0,io_cin[21]}; // @[Cat.scala 30:58]
  wire  ly6_out = ly6_in[0] ^ ly6_in[1] ^ ly6_in[2]; // @[CNN_CONV.scala 59:11]
  wire  out_cout_23 = ly6_in[0] & ly6_in[1] | ly6_in[0] & ly6_in[2] | ly6_in[1] & ly6_in[2]; // @[CNN_CONV.scala 64:21]
  wire [2:0] ly7_in = {ly6_out,io_cin[23:22]}; // @[Cat.scala 30:58]
  wire [9:0] _T_345 = {out_cout_9,out_cout_8,out_cout_7,out_cout_6,out_cout_5,out_cout_4,out_cout_3,out_cout_2,
    out_cout_1,out_cout_0}; // @[Cat.scala 30:58]
  wire [18:0] _T_354 = {out_cout_18,out_cout_17,out_cout_16,out_cout_15,out_cout_14,out_cout_13,out_cout_12,out_cout_11,
    out_cout_10,_T_345}; // @[Cat.scala 30:58]
  wire [22:0] _T_358 = {out_cout_22,out_cout_21,out_cout_20,out_cout_19,_T_354}; // @[Cat.scala 30:58]
  assign io_s = ly7_in[0] ^ ly7_in[1] ^ ly7_in[2]; // @[CNN_CONV.scala 59:11]
  assign io_c = ly7_in[0] & ly7_in[1] | ly7_in[0] & ly7_in[2] | ly7_in[1] & ly7_in[2]; // @[CNN_CONV.scala 64:21]
  assign io_cout = {out_cout_23,_T_358}; // @[Cat.scala 30:58]
endmodule
module WallaceAdder(
  input  [31:0] io_data_0,
  input  [31:0] io_data_1,
  input  [31:0] io_data_2,
  input  [31:0] io_data_3,
  input  [31:0] io_data_4,
  input  [31:0] io_data_5,
  input  [31:0] io_data_6,
  input  [31:0] io_data_7,
  input  [31:0] io_data_8,
  input  [31:0] io_data_9,
  input  [31:0] io_data_10,
  input  [31:0] io_data_11,
  input  [31:0] io_data_12,
  input  [31:0] io_data_13,
  input  [31:0] io_data_14,
  input  [31:0] io_data_15,
  input  [31:0] io_data_16,
  input  [31:0] io_data_17,
  input  [31:0] io_data_18,
  input  [31:0] io_data_19,
  input  [31:0] io_data_20,
  input  [31:0] io_data_21,
  input  [31:0] io_data_22,
  input  [31:0] io_data_23,
  input  [31:0] io_data_24,
  input         io_cin_0,
  input         io_cin_1,
  input         io_cin_2,
  input         io_cin_3,
  input         io_cin_4,
  input         io_cin_5,
  input         io_cin_6,
  input         io_cin_7,
  input         io_cin_8,
  input         io_cin_9,
  input         io_cin_10,
  input         io_cin_11,
  input         io_cin_12,
  input         io_cin_13,
  input         io_cin_14,
  input         io_cin_15,
  input         io_cin_16,
  input         io_cin_17,
  input         io_cin_18,
  input         io_cin_19,
  input         io_cin_20,
  input         io_cin_21,
  input         io_cin_22,
  input         io_cin_23,
  input         io_cin_24,
  output [31:0] io_s,
  output [31:0] io_c
);
  wire [24:0] WallaceTree25_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_1_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_1_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_1_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_1_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_1_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_2_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_2_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_2_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_2_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_2_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_3_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_3_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_3_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_3_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_3_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_4_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_4_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_4_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_4_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_4_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_5_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_5_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_5_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_5_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_5_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_6_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_6_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_6_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_6_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_6_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_7_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_7_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_7_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_7_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_7_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_8_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_8_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_8_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_8_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_8_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_9_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_9_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_9_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_9_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_9_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_10_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_10_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_10_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_10_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_10_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_11_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_11_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_11_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_11_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_11_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_12_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_12_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_12_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_12_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_12_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_13_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_13_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_13_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_13_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_13_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_14_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_14_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_14_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_14_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_14_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_15_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_15_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_15_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_15_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_15_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_16_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_16_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_16_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_16_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_16_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_17_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_17_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_17_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_17_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_17_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_18_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_18_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_18_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_18_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_18_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_19_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_19_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_19_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_19_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_19_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_20_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_20_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_20_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_20_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_20_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_21_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_21_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_21_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_21_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_21_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_22_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_22_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_22_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_22_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_22_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_23_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_23_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_23_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_23_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_23_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_24_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_24_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_24_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_24_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_24_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_25_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_25_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_25_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_25_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_25_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_26_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_26_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_26_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_26_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_26_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_27_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_27_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_27_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_27_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_27_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_28_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_28_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_28_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_28_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_28_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_29_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_29_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_29_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_29_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_29_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_30_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_30_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_30_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_30_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_30_io_cout; // @[CNN_CONV.scala 161:49]
  wire [24:0] WallaceTree25_31_io_n; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_31_io_cin; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_31_io_s; // @[CNN_CONV.scala 161:49]
  wire  WallaceTree25_31_io_c; // @[CNN_CONV.scala 161:49]
  wire [23:0] WallaceTree25_31_io_cout; // @[CNN_CONV.scala 161:49]
  wire [9:0] _T_8 = {io_cin_9,io_cin_8,io_cin_7,io_cin_6,io_cin_5,io_cin_4,io_cin_3,io_cin_2,io_cin_1,io_cin_0}; // @[Cat.scala 30:58]
  wire [18:0] _T_17 = {io_cin_18,io_cin_17,io_cin_16,io_cin_15,io_cin_14,io_cin_13,io_cin_12,io_cin_11,io_cin_10,_T_8}; // @[Cat.scala 30:58]
  wire [24:0] _T_23 = {io_cin_24,io_cin_23,io_cin_22,io_cin_21,io_cin_20,io_cin_19,_T_17}; // @[Cat.scala 30:58]
  wire [9:0] _T_58 = {io_data_9[0],io_data_8[0],io_data_7[0],io_data_6[0],io_data_5[0],io_data_4[0],io_data_3[0],
    io_data_2[0],io_data_1[0],io_data_0[0]}; // @[Cat.scala 30:58]
  wire [18:0] _T_67 = {io_data_18[0],io_data_17[0],io_data_16[0],io_data_15[0],io_data_14[0],io_data_13[0],io_data_12[0]
    ,io_data_11[0],io_data_10[0],_T_58}; // @[Cat.scala 30:58]
  wire [23:0] _T_72 = {io_data_23[0],io_data_22[0],io_data_21[0],io_data_20[0],io_data_19[0],_T_67}; // @[Cat.scala 30:58]
  wire [9:0] _T_107 = {io_data_9[1],io_data_8[1],io_data_7[1],io_data_6[1],io_data_5[1],io_data_4[1],io_data_3[1],
    io_data_2[1],io_data_1[1],io_data_0[1]}; // @[Cat.scala 30:58]
  wire [18:0] _T_116 = {io_data_18[1],io_data_17[1],io_data_16[1],io_data_15[1],io_data_14[1],io_data_13[1],io_data_12[1
    ],io_data_11[1],io_data_10[1],_T_107}; // @[Cat.scala 30:58]
  wire [23:0] _T_121 = {io_data_23[1],io_data_22[1],io_data_21[1],io_data_20[1],io_data_19[1],_T_116}; // @[Cat.scala 30:58]
  wire [9:0] _T_156 = {io_data_9[2],io_data_8[2],io_data_7[2],io_data_6[2],io_data_5[2],io_data_4[2],io_data_3[2],
    io_data_2[2],io_data_1[2],io_data_0[2]}; // @[Cat.scala 30:58]
  wire [18:0] _T_165 = {io_data_18[2],io_data_17[2],io_data_16[2],io_data_15[2],io_data_14[2],io_data_13[2],io_data_12[2
    ],io_data_11[2],io_data_10[2],_T_156}; // @[Cat.scala 30:58]
  wire [23:0] _T_170 = {io_data_23[2],io_data_22[2],io_data_21[2],io_data_20[2],io_data_19[2],_T_165}; // @[Cat.scala 30:58]
  wire [9:0] _T_205 = {io_data_9[3],io_data_8[3],io_data_7[3],io_data_6[3],io_data_5[3],io_data_4[3],io_data_3[3],
    io_data_2[3],io_data_1[3],io_data_0[3]}; // @[Cat.scala 30:58]
  wire [18:0] _T_214 = {io_data_18[3],io_data_17[3],io_data_16[3],io_data_15[3],io_data_14[3],io_data_13[3],io_data_12[3
    ],io_data_11[3],io_data_10[3],_T_205}; // @[Cat.scala 30:58]
  wire [23:0] _T_219 = {io_data_23[3],io_data_22[3],io_data_21[3],io_data_20[3],io_data_19[3],_T_214}; // @[Cat.scala 30:58]
  wire [9:0] _T_254 = {io_data_9[4],io_data_8[4],io_data_7[4],io_data_6[4],io_data_5[4],io_data_4[4],io_data_3[4],
    io_data_2[4],io_data_1[4],io_data_0[4]}; // @[Cat.scala 30:58]
  wire [18:0] _T_263 = {io_data_18[4],io_data_17[4],io_data_16[4],io_data_15[4],io_data_14[4],io_data_13[4],io_data_12[4
    ],io_data_11[4],io_data_10[4],_T_254}; // @[Cat.scala 30:58]
  wire [23:0] _T_268 = {io_data_23[4],io_data_22[4],io_data_21[4],io_data_20[4],io_data_19[4],_T_263}; // @[Cat.scala 30:58]
  wire [9:0] _T_303 = {io_data_9[5],io_data_8[5],io_data_7[5],io_data_6[5],io_data_5[5],io_data_4[5],io_data_3[5],
    io_data_2[5],io_data_1[5],io_data_0[5]}; // @[Cat.scala 30:58]
  wire [18:0] _T_312 = {io_data_18[5],io_data_17[5],io_data_16[5],io_data_15[5],io_data_14[5],io_data_13[5],io_data_12[5
    ],io_data_11[5],io_data_10[5],_T_303}; // @[Cat.scala 30:58]
  wire [23:0] _T_317 = {io_data_23[5],io_data_22[5],io_data_21[5],io_data_20[5],io_data_19[5],_T_312}; // @[Cat.scala 30:58]
  wire [9:0] _T_352 = {io_data_9[6],io_data_8[6],io_data_7[6],io_data_6[6],io_data_5[6],io_data_4[6],io_data_3[6],
    io_data_2[6],io_data_1[6],io_data_0[6]}; // @[Cat.scala 30:58]
  wire [18:0] _T_361 = {io_data_18[6],io_data_17[6],io_data_16[6],io_data_15[6],io_data_14[6],io_data_13[6],io_data_12[6
    ],io_data_11[6],io_data_10[6],_T_352}; // @[Cat.scala 30:58]
  wire [23:0] _T_366 = {io_data_23[6],io_data_22[6],io_data_21[6],io_data_20[6],io_data_19[6],_T_361}; // @[Cat.scala 30:58]
  wire [9:0] _T_401 = {io_data_9[7],io_data_8[7],io_data_7[7],io_data_6[7],io_data_5[7],io_data_4[7],io_data_3[7],
    io_data_2[7],io_data_1[7],io_data_0[7]}; // @[Cat.scala 30:58]
  wire [18:0] _T_410 = {io_data_18[7],io_data_17[7],io_data_16[7],io_data_15[7],io_data_14[7],io_data_13[7],io_data_12[7
    ],io_data_11[7],io_data_10[7],_T_401}; // @[Cat.scala 30:58]
  wire [23:0] _T_415 = {io_data_23[7],io_data_22[7],io_data_21[7],io_data_20[7],io_data_19[7],_T_410}; // @[Cat.scala 30:58]
  wire [9:0] _T_450 = {io_data_9[8],io_data_8[8],io_data_7[8],io_data_6[8],io_data_5[8],io_data_4[8],io_data_3[8],
    io_data_2[8],io_data_1[8],io_data_0[8]}; // @[Cat.scala 30:58]
  wire [18:0] _T_459 = {io_data_18[8],io_data_17[8],io_data_16[8],io_data_15[8],io_data_14[8],io_data_13[8],io_data_12[8
    ],io_data_11[8],io_data_10[8],_T_450}; // @[Cat.scala 30:58]
  wire [23:0] _T_464 = {io_data_23[8],io_data_22[8],io_data_21[8],io_data_20[8],io_data_19[8],_T_459}; // @[Cat.scala 30:58]
  wire [9:0] _T_499 = {io_data_9[9],io_data_8[9],io_data_7[9],io_data_6[9],io_data_5[9],io_data_4[9],io_data_3[9],
    io_data_2[9],io_data_1[9],io_data_0[9]}; // @[Cat.scala 30:58]
  wire [18:0] _T_508 = {io_data_18[9],io_data_17[9],io_data_16[9],io_data_15[9],io_data_14[9],io_data_13[9],io_data_12[9
    ],io_data_11[9],io_data_10[9],_T_499}; // @[Cat.scala 30:58]
  wire [23:0] _T_513 = {io_data_23[9],io_data_22[9],io_data_21[9],io_data_20[9],io_data_19[9],_T_508}; // @[Cat.scala 30:58]
  wire [9:0] _T_548 = {io_data_9[10],io_data_8[10],io_data_7[10],io_data_6[10],io_data_5[10],io_data_4[10],io_data_3[10]
    ,io_data_2[10],io_data_1[10],io_data_0[10]}; // @[Cat.scala 30:58]
  wire [18:0] _T_557 = {io_data_18[10],io_data_17[10],io_data_16[10],io_data_15[10],io_data_14[10],io_data_13[10],
    io_data_12[10],io_data_11[10],io_data_10[10],_T_548}; // @[Cat.scala 30:58]
  wire [23:0] _T_562 = {io_data_23[10],io_data_22[10],io_data_21[10],io_data_20[10],io_data_19[10],_T_557}; // @[Cat.scala 30:58]
  wire [9:0] _T_597 = {io_data_9[11],io_data_8[11],io_data_7[11],io_data_6[11],io_data_5[11],io_data_4[11],io_data_3[11]
    ,io_data_2[11],io_data_1[11],io_data_0[11]}; // @[Cat.scala 30:58]
  wire [18:0] _T_606 = {io_data_18[11],io_data_17[11],io_data_16[11],io_data_15[11],io_data_14[11],io_data_13[11],
    io_data_12[11],io_data_11[11],io_data_10[11],_T_597}; // @[Cat.scala 30:58]
  wire [23:0] _T_611 = {io_data_23[11],io_data_22[11],io_data_21[11],io_data_20[11],io_data_19[11],_T_606}; // @[Cat.scala 30:58]
  wire [9:0] _T_646 = {io_data_9[12],io_data_8[12],io_data_7[12],io_data_6[12],io_data_5[12],io_data_4[12],io_data_3[12]
    ,io_data_2[12],io_data_1[12],io_data_0[12]}; // @[Cat.scala 30:58]
  wire [18:0] _T_655 = {io_data_18[12],io_data_17[12],io_data_16[12],io_data_15[12],io_data_14[12],io_data_13[12],
    io_data_12[12],io_data_11[12],io_data_10[12],_T_646}; // @[Cat.scala 30:58]
  wire [23:0] _T_660 = {io_data_23[12],io_data_22[12],io_data_21[12],io_data_20[12],io_data_19[12],_T_655}; // @[Cat.scala 30:58]
  wire [9:0] _T_695 = {io_data_9[13],io_data_8[13],io_data_7[13],io_data_6[13],io_data_5[13],io_data_4[13],io_data_3[13]
    ,io_data_2[13],io_data_1[13],io_data_0[13]}; // @[Cat.scala 30:58]
  wire [18:0] _T_704 = {io_data_18[13],io_data_17[13],io_data_16[13],io_data_15[13],io_data_14[13],io_data_13[13],
    io_data_12[13],io_data_11[13],io_data_10[13],_T_695}; // @[Cat.scala 30:58]
  wire [23:0] _T_709 = {io_data_23[13],io_data_22[13],io_data_21[13],io_data_20[13],io_data_19[13],_T_704}; // @[Cat.scala 30:58]
  wire [9:0] _T_744 = {io_data_9[14],io_data_8[14],io_data_7[14],io_data_6[14],io_data_5[14],io_data_4[14],io_data_3[14]
    ,io_data_2[14],io_data_1[14],io_data_0[14]}; // @[Cat.scala 30:58]
  wire [18:0] _T_753 = {io_data_18[14],io_data_17[14],io_data_16[14],io_data_15[14],io_data_14[14],io_data_13[14],
    io_data_12[14],io_data_11[14],io_data_10[14],_T_744}; // @[Cat.scala 30:58]
  wire [23:0] _T_758 = {io_data_23[14],io_data_22[14],io_data_21[14],io_data_20[14],io_data_19[14],_T_753}; // @[Cat.scala 30:58]
  wire [9:0] _T_793 = {io_data_9[15],io_data_8[15],io_data_7[15],io_data_6[15],io_data_5[15],io_data_4[15],io_data_3[15]
    ,io_data_2[15],io_data_1[15],io_data_0[15]}; // @[Cat.scala 30:58]
  wire [18:0] _T_802 = {io_data_18[15],io_data_17[15],io_data_16[15],io_data_15[15],io_data_14[15],io_data_13[15],
    io_data_12[15],io_data_11[15],io_data_10[15],_T_793}; // @[Cat.scala 30:58]
  wire [23:0] _T_807 = {io_data_23[15],io_data_22[15],io_data_21[15],io_data_20[15],io_data_19[15],_T_802}; // @[Cat.scala 30:58]
  wire [9:0] _T_842 = {io_data_9[16],io_data_8[16],io_data_7[16],io_data_6[16],io_data_5[16],io_data_4[16],io_data_3[16]
    ,io_data_2[16],io_data_1[16],io_data_0[16]}; // @[Cat.scala 30:58]
  wire [18:0] _T_851 = {io_data_18[16],io_data_17[16],io_data_16[16],io_data_15[16],io_data_14[16],io_data_13[16],
    io_data_12[16],io_data_11[16],io_data_10[16],_T_842}; // @[Cat.scala 30:58]
  wire [23:0] _T_856 = {io_data_23[16],io_data_22[16],io_data_21[16],io_data_20[16],io_data_19[16],_T_851}; // @[Cat.scala 30:58]
  wire [9:0] _T_891 = {io_data_9[17],io_data_8[17],io_data_7[17],io_data_6[17],io_data_5[17],io_data_4[17],io_data_3[17]
    ,io_data_2[17],io_data_1[17],io_data_0[17]}; // @[Cat.scala 30:58]
  wire [18:0] _T_900 = {io_data_18[17],io_data_17[17],io_data_16[17],io_data_15[17],io_data_14[17],io_data_13[17],
    io_data_12[17],io_data_11[17],io_data_10[17],_T_891}; // @[Cat.scala 30:58]
  wire [23:0] _T_905 = {io_data_23[17],io_data_22[17],io_data_21[17],io_data_20[17],io_data_19[17],_T_900}; // @[Cat.scala 30:58]
  wire [9:0] _T_940 = {io_data_9[18],io_data_8[18],io_data_7[18],io_data_6[18],io_data_5[18],io_data_4[18],io_data_3[18]
    ,io_data_2[18],io_data_1[18],io_data_0[18]}; // @[Cat.scala 30:58]
  wire [18:0] _T_949 = {io_data_18[18],io_data_17[18],io_data_16[18],io_data_15[18],io_data_14[18],io_data_13[18],
    io_data_12[18],io_data_11[18],io_data_10[18],_T_940}; // @[Cat.scala 30:58]
  wire [23:0] _T_954 = {io_data_23[18],io_data_22[18],io_data_21[18],io_data_20[18],io_data_19[18],_T_949}; // @[Cat.scala 30:58]
  wire [9:0] _T_989 = {io_data_9[19],io_data_8[19],io_data_7[19],io_data_6[19],io_data_5[19],io_data_4[19],io_data_3[19]
    ,io_data_2[19],io_data_1[19],io_data_0[19]}; // @[Cat.scala 30:58]
  wire [18:0] _T_998 = {io_data_18[19],io_data_17[19],io_data_16[19],io_data_15[19],io_data_14[19],io_data_13[19],
    io_data_12[19],io_data_11[19],io_data_10[19],_T_989}; // @[Cat.scala 30:58]
  wire [23:0] _T_1003 = {io_data_23[19],io_data_22[19],io_data_21[19],io_data_20[19],io_data_19[19],_T_998}; // @[Cat.scala 30:58]
  wire [9:0] _T_1038 = {io_data_9[20],io_data_8[20],io_data_7[20],io_data_6[20],io_data_5[20],io_data_4[20],io_data_3[20
    ],io_data_2[20],io_data_1[20],io_data_0[20]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1047 = {io_data_18[20],io_data_17[20],io_data_16[20],io_data_15[20],io_data_14[20],io_data_13[20],
    io_data_12[20],io_data_11[20],io_data_10[20],_T_1038}; // @[Cat.scala 30:58]
  wire [23:0] _T_1052 = {io_data_23[20],io_data_22[20],io_data_21[20],io_data_20[20],io_data_19[20],_T_1047}; // @[Cat.scala 30:58]
  wire [9:0] _T_1087 = {io_data_9[21],io_data_8[21],io_data_7[21],io_data_6[21],io_data_5[21],io_data_4[21],io_data_3[21
    ],io_data_2[21],io_data_1[21],io_data_0[21]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1096 = {io_data_18[21],io_data_17[21],io_data_16[21],io_data_15[21],io_data_14[21],io_data_13[21],
    io_data_12[21],io_data_11[21],io_data_10[21],_T_1087}; // @[Cat.scala 30:58]
  wire [23:0] _T_1101 = {io_data_23[21],io_data_22[21],io_data_21[21],io_data_20[21],io_data_19[21],_T_1096}; // @[Cat.scala 30:58]
  wire [9:0] _T_1136 = {io_data_9[22],io_data_8[22],io_data_7[22],io_data_6[22],io_data_5[22],io_data_4[22],io_data_3[22
    ],io_data_2[22],io_data_1[22],io_data_0[22]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1145 = {io_data_18[22],io_data_17[22],io_data_16[22],io_data_15[22],io_data_14[22],io_data_13[22],
    io_data_12[22],io_data_11[22],io_data_10[22],_T_1136}; // @[Cat.scala 30:58]
  wire [23:0] _T_1150 = {io_data_23[22],io_data_22[22],io_data_21[22],io_data_20[22],io_data_19[22],_T_1145}; // @[Cat.scala 30:58]
  wire [9:0] _T_1185 = {io_data_9[23],io_data_8[23],io_data_7[23],io_data_6[23],io_data_5[23],io_data_4[23],io_data_3[23
    ],io_data_2[23],io_data_1[23],io_data_0[23]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1194 = {io_data_18[23],io_data_17[23],io_data_16[23],io_data_15[23],io_data_14[23],io_data_13[23],
    io_data_12[23],io_data_11[23],io_data_10[23],_T_1185}; // @[Cat.scala 30:58]
  wire [23:0] _T_1199 = {io_data_23[23],io_data_22[23],io_data_21[23],io_data_20[23],io_data_19[23],_T_1194}; // @[Cat.scala 30:58]
  wire [9:0] _T_1234 = {io_data_9[24],io_data_8[24],io_data_7[24],io_data_6[24],io_data_5[24],io_data_4[24],io_data_3[24
    ],io_data_2[24],io_data_1[24],io_data_0[24]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1243 = {io_data_18[24],io_data_17[24],io_data_16[24],io_data_15[24],io_data_14[24],io_data_13[24],
    io_data_12[24],io_data_11[24],io_data_10[24],_T_1234}; // @[Cat.scala 30:58]
  wire [23:0] _T_1248 = {io_data_23[24],io_data_22[24],io_data_21[24],io_data_20[24],io_data_19[24],_T_1243}; // @[Cat.scala 30:58]
  wire [9:0] _T_1283 = {io_data_9[25],io_data_8[25],io_data_7[25],io_data_6[25],io_data_5[25],io_data_4[25],io_data_3[25
    ],io_data_2[25],io_data_1[25],io_data_0[25]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1292 = {io_data_18[25],io_data_17[25],io_data_16[25],io_data_15[25],io_data_14[25],io_data_13[25],
    io_data_12[25],io_data_11[25],io_data_10[25],_T_1283}; // @[Cat.scala 30:58]
  wire [23:0] _T_1297 = {io_data_23[25],io_data_22[25],io_data_21[25],io_data_20[25],io_data_19[25],_T_1292}; // @[Cat.scala 30:58]
  wire [9:0] _T_1332 = {io_data_9[26],io_data_8[26],io_data_7[26],io_data_6[26],io_data_5[26],io_data_4[26],io_data_3[26
    ],io_data_2[26],io_data_1[26],io_data_0[26]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1341 = {io_data_18[26],io_data_17[26],io_data_16[26],io_data_15[26],io_data_14[26],io_data_13[26],
    io_data_12[26],io_data_11[26],io_data_10[26],_T_1332}; // @[Cat.scala 30:58]
  wire [23:0] _T_1346 = {io_data_23[26],io_data_22[26],io_data_21[26],io_data_20[26],io_data_19[26],_T_1341}; // @[Cat.scala 30:58]
  wire [9:0] _T_1381 = {io_data_9[27],io_data_8[27],io_data_7[27],io_data_6[27],io_data_5[27],io_data_4[27],io_data_3[27
    ],io_data_2[27],io_data_1[27],io_data_0[27]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1390 = {io_data_18[27],io_data_17[27],io_data_16[27],io_data_15[27],io_data_14[27],io_data_13[27],
    io_data_12[27],io_data_11[27],io_data_10[27],_T_1381}; // @[Cat.scala 30:58]
  wire [23:0] _T_1395 = {io_data_23[27],io_data_22[27],io_data_21[27],io_data_20[27],io_data_19[27],_T_1390}; // @[Cat.scala 30:58]
  wire [9:0] _T_1430 = {io_data_9[28],io_data_8[28],io_data_7[28],io_data_6[28],io_data_5[28],io_data_4[28],io_data_3[28
    ],io_data_2[28],io_data_1[28],io_data_0[28]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1439 = {io_data_18[28],io_data_17[28],io_data_16[28],io_data_15[28],io_data_14[28],io_data_13[28],
    io_data_12[28],io_data_11[28],io_data_10[28],_T_1430}; // @[Cat.scala 30:58]
  wire [23:0] _T_1444 = {io_data_23[28],io_data_22[28],io_data_21[28],io_data_20[28],io_data_19[28],_T_1439}; // @[Cat.scala 30:58]
  wire [9:0] _T_1479 = {io_data_9[29],io_data_8[29],io_data_7[29],io_data_6[29],io_data_5[29],io_data_4[29],io_data_3[29
    ],io_data_2[29],io_data_1[29],io_data_0[29]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1488 = {io_data_18[29],io_data_17[29],io_data_16[29],io_data_15[29],io_data_14[29],io_data_13[29],
    io_data_12[29],io_data_11[29],io_data_10[29],_T_1479}; // @[Cat.scala 30:58]
  wire [23:0] _T_1493 = {io_data_23[29],io_data_22[29],io_data_21[29],io_data_20[29],io_data_19[29],_T_1488}; // @[Cat.scala 30:58]
  wire [9:0] _T_1528 = {io_data_9[30],io_data_8[30],io_data_7[30],io_data_6[30],io_data_5[30],io_data_4[30],io_data_3[30
    ],io_data_2[30],io_data_1[30],io_data_0[30]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1537 = {io_data_18[30],io_data_17[30],io_data_16[30],io_data_15[30],io_data_14[30],io_data_13[30],
    io_data_12[30],io_data_11[30],io_data_10[30],_T_1528}; // @[Cat.scala 30:58]
  wire [23:0] _T_1542 = {io_data_23[30],io_data_22[30],io_data_21[30],io_data_20[30],io_data_19[30],_T_1537}; // @[Cat.scala 30:58]
  wire [9:0] _T_1577 = {io_data_9[31],io_data_8[31],io_data_7[31],io_data_6[31],io_data_5[31],io_data_4[31],io_data_3[31
    ],io_data_2[31],io_data_1[31],io_data_0[31]}; // @[Cat.scala 30:58]
  wire [18:0] _T_1586 = {io_data_18[31],io_data_17[31],io_data_16[31],io_data_15[31],io_data_14[31],io_data_13[31],
    io_data_12[31],io_data_11[31],io_data_10[31],_T_1577}; // @[Cat.scala 30:58]
  wire [23:0] _T_1591 = {io_data_23[31],io_data_22[31],io_data_21[31],io_data_20[31],io_data_19[31],_T_1586}; // @[Cat.scala 30:58]
  wire  wallace_tree_1_s = WallaceTree25_1_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_0_s = WallaceTree25_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_2_s = WallaceTree25_2_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_3_s = WallaceTree25_3_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_4_s = WallaceTree25_4_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_5_s = WallaceTree25_5_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_6_s = WallaceTree25_6_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_7_s = WallaceTree25_7_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_8_s = WallaceTree25_8_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_9_s = WallaceTree25_9_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire [9:0] _T_1601 = {wallace_tree_9_s,wallace_tree_8_s,wallace_tree_7_s,wallace_tree_6_s,wallace_tree_5_s,
    wallace_tree_4_s,wallace_tree_3_s,wallace_tree_2_s,wallace_tree_1_s,wallace_tree_0_s}; // @[Cat.scala 30:58]
  wire  wallace_tree_10_s = WallaceTree25_10_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_11_s = WallaceTree25_11_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_12_s = WallaceTree25_12_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_13_s = WallaceTree25_13_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_14_s = WallaceTree25_14_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_15_s = WallaceTree25_15_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_16_s = WallaceTree25_16_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_17_s = WallaceTree25_17_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_18_s = WallaceTree25_18_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire [18:0] _T_1610 = {wallace_tree_18_s,wallace_tree_17_s,wallace_tree_16_s,wallace_tree_15_s,wallace_tree_14_s,
    wallace_tree_13_s,wallace_tree_12_s,wallace_tree_11_s,wallace_tree_10_s,_T_1601}; // @[Cat.scala 30:58]
  wire  wallace_tree_19_s = WallaceTree25_19_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_20_s = WallaceTree25_20_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_21_s = WallaceTree25_21_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_22_s = WallaceTree25_22_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_23_s = WallaceTree25_23_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_24_s = WallaceTree25_24_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_25_s = WallaceTree25_25_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_26_s = WallaceTree25_26_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_27_s = WallaceTree25_27_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire [27:0] _T_1619 = {wallace_tree_27_s,wallace_tree_26_s,wallace_tree_25_s,wallace_tree_24_s,wallace_tree_23_s,
    wallace_tree_22_s,wallace_tree_21_s,wallace_tree_20_s,wallace_tree_19_s,_T_1610}; // @[Cat.scala 30:58]
  wire  wallace_tree_28_s = WallaceTree25_28_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_29_s = WallaceTree25_29_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_30_s = WallaceTree25_30_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire [30:0] _T_1622 = {wallace_tree_30_s,wallace_tree_29_s,wallace_tree_28_s,_T_1619}; // @[Cat.scala 30:58]
  wire  wallace_tree_31_s = WallaceTree25_31_io_s; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_0_c = WallaceTree25_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_1_c = WallaceTree25_1_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_2_c = WallaceTree25_2_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_3_c = WallaceTree25_3_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_4_c = WallaceTree25_4_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_5_c = WallaceTree25_5_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_6_c = WallaceTree25_6_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_7_c = WallaceTree25_7_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_8_c = WallaceTree25_8_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire [9:0] _T_1632 = {wallace_tree_8_c,wallace_tree_7_c,wallace_tree_6_c,wallace_tree_5_c,wallace_tree_4_c,
    wallace_tree_3_c,wallace_tree_2_c,wallace_tree_1_c,wallace_tree_0_c,io_cin_24}; // @[Cat.scala 30:58]
  wire  wallace_tree_9_c = WallaceTree25_9_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_10_c = WallaceTree25_10_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_11_c = WallaceTree25_11_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_12_c = WallaceTree25_12_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_13_c = WallaceTree25_13_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_14_c = WallaceTree25_14_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_15_c = WallaceTree25_15_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_16_c = WallaceTree25_16_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_17_c = WallaceTree25_17_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire [18:0] _T_1641 = {wallace_tree_17_c,wallace_tree_16_c,wallace_tree_15_c,wallace_tree_14_c,wallace_tree_13_c,
    wallace_tree_12_c,wallace_tree_11_c,wallace_tree_10_c,wallace_tree_9_c,_T_1632}; // @[Cat.scala 30:58]
  wire  wallace_tree_18_c = WallaceTree25_18_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_19_c = WallaceTree25_19_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_20_c = WallaceTree25_20_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_21_c = WallaceTree25_21_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_22_c = WallaceTree25_22_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_23_c = WallaceTree25_23_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_24_c = WallaceTree25_24_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_25_c = WallaceTree25_25_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_26_c = WallaceTree25_26_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire [27:0] _T_1650 = {wallace_tree_26_c,wallace_tree_25_c,wallace_tree_24_c,wallace_tree_23_c,wallace_tree_22_c,
    wallace_tree_21_c,wallace_tree_20_c,wallace_tree_19_c,wallace_tree_18_c,_T_1641}; // @[Cat.scala 30:58]
  wire  wallace_tree_27_c = WallaceTree25_27_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_28_c = WallaceTree25_28_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire  wallace_tree_29_c = WallaceTree25_29_io_c; // @[CNN_CONV.scala 161:{29,29}]
  wire [30:0] _T_1653 = {wallace_tree_29_c,wallace_tree_28_c,wallace_tree_27_c,_T_1650}; // @[Cat.scala 30:58]
  wire  wallace_tree_30_c = WallaceTree25_30_io_c; // @[CNN_CONV.scala 161:{29,29}]
  WallaceTree25 WallaceTree25 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_io_n),
    .io_cin(WallaceTree25_io_cin),
    .io_s(WallaceTree25_io_s),
    .io_c(WallaceTree25_io_c),
    .io_cout(WallaceTree25_io_cout)
  );
  WallaceTree25 WallaceTree25_1 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_1_io_n),
    .io_cin(WallaceTree25_1_io_cin),
    .io_s(WallaceTree25_1_io_s),
    .io_c(WallaceTree25_1_io_c),
    .io_cout(WallaceTree25_1_io_cout)
  );
  WallaceTree25 WallaceTree25_2 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_2_io_n),
    .io_cin(WallaceTree25_2_io_cin),
    .io_s(WallaceTree25_2_io_s),
    .io_c(WallaceTree25_2_io_c),
    .io_cout(WallaceTree25_2_io_cout)
  );
  WallaceTree25 WallaceTree25_3 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_3_io_n),
    .io_cin(WallaceTree25_3_io_cin),
    .io_s(WallaceTree25_3_io_s),
    .io_c(WallaceTree25_3_io_c),
    .io_cout(WallaceTree25_3_io_cout)
  );
  WallaceTree25 WallaceTree25_4 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_4_io_n),
    .io_cin(WallaceTree25_4_io_cin),
    .io_s(WallaceTree25_4_io_s),
    .io_c(WallaceTree25_4_io_c),
    .io_cout(WallaceTree25_4_io_cout)
  );
  WallaceTree25 WallaceTree25_5 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_5_io_n),
    .io_cin(WallaceTree25_5_io_cin),
    .io_s(WallaceTree25_5_io_s),
    .io_c(WallaceTree25_5_io_c),
    .io_cout(WallaceTree25_5_io_cout)
  );
  WallaceTree25 WallaceTree25_6 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_6_io_n),
    .io_cin(WallaceTree25_6_io_cin),
    .io_s(WallaceTree25_6_io_s),
    .io_c(WallaceTree25_6_io_c),
    .io_cout(WallaceTree25_6_io_cout)
  );
  WallaceTree25 WallaceTree25_7 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_7_io_n),
    .io_cin(WallaceTree25_7_io_cin),
    .io_s(WallaceTree25_7_io_s),
    .io_c(WallaceTree25_7_io_c),
    .io_cout(WallaceTree25_7_io_cout)
  );
  WallaceTree25 WallaceTree25_8 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_8_io_n),
    .io_cin(WallaceTree25_8_io_cin),
    .io_s(WallaceTree25_8_io_s),
    .io_c(WallaceTree25_8_io_c),
    .io_cout(WallaceTree25_8_io_cout)
  );
  WallaceTree25 WallaceTree25_9 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_9_io_n),
    .io_cin(WallaceTree25_9_io_cin),
    .io_s(WallaceTree25_9_io_s),
    .io_c(WallaceTree25_9_io_c),
    .io_cout(WallaceTree25_9_io_cout)
  );
  WallaceTree25 WallaceTree25_10 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_10_io_n),
    .io_cin(WallaceTree25_10_io_cin),
    .io_s(WallaceTree25_10_io_s),
    .io_c(WallaceTree25_10_io_c),
    .io_cout(WallaceTree25_10_io_cout)
  );
  WallaceTree25 WallaceTree25_11 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_11_io_n),
    .io_cin(WallaceTree25_11_io_cin),
    .io_s(WallaceTree25_11_io_s),
    .io_c(WallaceTree25_11_io_c),
    .io_cout(WallaceTree25_11_io_cout)
  );
  WallaceTree25 WallaceTree25_12 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_12_io_n),
    .io_cin(WallaceTree25_12_io_cin),
    .io_s(WallaceTree25_12_io_s),
    .io_c(WallaceTree25_12_io_c),
    .io_cout(WallaceTree25_12_io_cout)
  );
  WallaceTree25 WallaceTree25_13 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_13_io_n),
    .io_cin(WallaceTree25_13_io_cin),
    .io_s(WallaceTree25_13_io_s),
    .io_c(WallaceTree25_13_io_c),
    .io_cout(WallaceTree25_13_io_cout)
  );
  WallaceTree25 WallaceTree25_14 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_14_io_n),
    .io_cin(WallaceTree25_14_io_cin),
    .io_s(WallaceTree25_14_io_s),
    .io_c(WallaceTree25_14_io_c),
    .io_cout(WallaceTree25_14_io_cout)
  );
  WallaceTree25 WallaceTree25_15 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_15_io_n),
    .io_cin(WallaceTree25_15_io_cin),
    .io_s(WallaceTree25_15_io_s),
    .io_c(WallaceTree25_15_io_c),
    .io_cout(WallaceTree25_15_io_cout)
  );
  WallaceTree25 WallaceTree25_16 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_16_io_n),
    .io_cin(WallaceTree25_16_io_cin),
    .io_s(WallaceTree25_16_io_s),
    .io_c(WallaceTree25_16_io_c),
    .io_cout(WallaceTree25_16_io_cout)
  );
  WallaceTree25 WallaceTree25_17 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_17_io_n),
    .io_cin(WallaceTree25_17_io_cin),
    .io_s(WallaceTree25_17_io_s),
    .io_c(WallaceTree25_17_io_c),
    .io_cout(WallaceTree25_17_io_cout)
  );
  WallaceTree25 WallaceTree25_18 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_18_io_n),
    .io_cin(WallaceTree25_18_io_cin),
    .io_s(WallaceTree25_18_io_s),
    .io_c(WallaceTree25_18_io_c),
    .io_cout(WallaceTree25_18_io_cout)
  );
  WallaceTree25 WallaceTree25_19 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_19_io_n),
    .io_cin(WallaceTree25_19_io_cin),
    .io_s(WallaceTree25_19_io_s),
    .io_c(WallaceTree25_19_io_c),
    .io_cout(WallaceTree25_19_io_cout)
  );
  WallaceTree25 WallaceTree25_20 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_20_io_n),
    .io_cin(WallaceTree25_20_io_cin),
    .io_s(WallaceTree25_20_io_s),
    .io_c(WallaceTree25_20_io_c),
    .io_cout(WallaceTree25_20_io_cout)
  );
  WallaceTree25 WallaceTree25_21 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_21_io_n),
    .io_cin(WallaceTree25_21_io_cin),
    .io_s(WallaceTree25_21_io_s),
    .io_c(WallaceTree25_21_io_c),
    .io_cout(WallaceTree25_21_io_cout)
  );
  WallaceTree25 WallaceTree25_22 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_22_io_n),
    .io_cin(WallaceTree25_22_io_cin),
    .io_s(WallaceTree25_22_io_s),
    .io_c(WallaceTree25_22_io_c),
    .io_cout(WallaceTree25_22_io_cout)
  );
  WallaceTree25 WallaceTree25_23 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_23_io_n),
    .io_cin(WallaceTree25_23_io_cin),
    .io_s(WallaceTree25_23_io_s),
    .io_c(WallaceTree25_23_io_c),
    .io_cout(WallaceTree25_23_io_cout)
  );
  WallaceTree25 WallaceTree25_24 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_24_io_n),
    .io_cin(WallaceTree25_24_io_cin),
    .io_s(WallaceTree25_24_io_s),
    .io_c(WallaceTree25_24_io_c),
    .io_cout(WallaceTree25_24_io_cout)
  );
  WallaceTree25 WallaceTree25_25 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_25_io_n),
    .io_cin(WallaceTree25_25_io_cin),
    .io_s(WallaceTree25_25_io_s),
    .io_c(WallaceTree25_25_io_c),
    .io_cout(WallaceTree25_25_io_cout)
  );
  WallaceTree25 WallaceTree25_26 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_26_io_n),
    .io_cin(WallaceTree25_26_io_cin),
    .io_s(WallaceTree25_26_io_s),
    .io_c(WallaceTree25_26_io_c),
    .io_cout(WallaceTree25_26_io_cout)
  );
  WallaceTree25 WallaceTree25_27 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_27_io_n),
    .io_cin(WallaceTree25_27_io_cin),
    .io_s(WallaceTree25_27_io_s),
    .io_c(WallaceTree25_27_io_c),
    .io_cout(WallaceTree25_27_io_cout)
  );
  WallaceTree25 WallaceTree25_28 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_28_io_n),
    .io_cin(WallaceTree25_28_io_cin),
    .io_s(WallaceTree25_28_io_s),
    .io_c(WallaceTree25_28_io_c),
    .io_cout(WallaceTree25_28_io_cout)
  );
  WallaceTree25 WallaceTree25_29 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_29_io_n),
    .io_cin(WallaceTree25_29_io_cin),
    .io_s(WallaceTree25_29_io_s),
    .io_c(WallaceTree25_29_io_c),
    .io_cout(WallaceTree25_29_io_cout)
  );
  WallaceTree25 WallaceTree25_30 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_30_io_n),
    .io_cin(WallaceTree25_30_io_cin),
    .io_s(WallaceTree25_30_io_s),
    .io_c(WallaceTree25_30_io_c),
    .io_cout(WallaceTree25_30_io_cout)
  );
  WallaceTree25 WallaceTree25_31 ( // @[CNN_CONV.scala 161:49]
    .io_n(WallaceTree25_31_io_n),
    .io_cin(WallaceTree25_31_io_cin),
    .io_s(WallaceTree25_31_io_s),
    .io_c(WallaceTree25_31_io_c),
    .io_cout(WallaceTree25_31_io_cout)
  );
  assign io_s = {wallace_tree_31_s,_T_1622}; // @[Cat.scala 30:58]
  assign io_c = {wallace_tree_30_c,_T_1653}; // @[Cat.scala 30:58]
  assign WallaceTree25_io_n = {io_data_24[0],_T_72}; // @[Cat.scala 30:58]
  assign WallaceTree25_io_cin = _T_23[23:0]; // @[CNN_CONV.scala 155:56]
  assign WallaceTree25_1_io_n = {io_data_24[1],_T_121}; // @[Cat.scala 30:58]
  assign WallaceTree25_1_io_cin = WallaceTree25_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_2_io_n = {io_data_24[2],_T_170}; // @[Cat.scala 30:58]
  assign WallaceTree25_2_io_cin = WallaceTree25_1_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_3_io_n = {io_data_24[3],_T_219}; // @[Cat.scala 30:58]
  assign WallaceTree25_3_io_cin = WallaceTree25_2_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_4_io_n = {io_data_24[4],_T_268}; // @[Cat.scala 30:58]
  assign WallaceTree25_4_io_cin = WallaceTree25_3_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_5_io_n = {io_data_24[5],_T_317}; // @[Cat.scala 30:58]
  assign WallaceTree25_5_io_cin = WallaceTree25_4_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_6_io_n = {io_data_24[6],_T_366}; // @[Cat.scala 30:58]
  assign WallaceTree25_6_io_cin = WallaceTree25_5_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_7_io_n = {io_data_24[7],_T_415}; // @[Cat.scala 30:58]
  assign WallaceTree25_7_io_cin = WallaceTree25_6_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_8_io_n = {io_data_24[8],_T_464}; // @[Cat.scala 30:58]
  assign WallaceTree25_8_io_cin = WallaceTree25_7_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_9_io_n = {io_data_24[9],_T_513}; // @[Cat.scala 30:58]
  assign WallaceTree25_9_io_cin = WallaceTree25_8_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_10_io_n = {io_data_24[10],_T_562}; // @[Cat.scala 30:58]
  assign WallaceTree25_10_io_cin = WallaceTree25_9_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_11_io_n = {io_data_24[11],_T_611}; // @[Cat.scala 30:58]
  assign WallaceTree25_11_io_cin = WallaceTree25_10_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_12_io_n = {io_data_24[12],_T_660}; // @[Cat.scala 30:58]
  assign WallaceTree25_12_io_cin = WallaceTree25_11_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_13_io_n = {io_data_24[13],_T_709}; // @[Cat.scala 30:58]
  assign WallaceTree25_13_io_cin = WallaceTree25_12_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_14_io_n = {io_data_24[14],_T_758}; // @[Cat.scala 30:58]
  assign WallaceTree25_14_io_cin = WallaceTree25_13_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_15_io_n = {io_data_24[15],_T_807}; // @[Cat.scala 30:58]
  assign WallaceTree25_15_io_cin = WallaceTree25_14_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_16_io_n = {io_data_24[16],_T_856}; // @[Cat.scala 30:58]
  assign WallaceTree25_16_io_cin = WallaceTree25_15_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_17_io_n = {io_data_24[17],_T_905}; // @[Cat.scala 30:58]
  assign WallaceTree25_17_io_cin = WallaceTree25_16_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_18_io_n = {io_data_24[18],_T_954}; // @[Cat.scala 30:58]
  assign WallaceTree25_18_io_cin = WallaceTree25_17_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_19_io_n = {io_data_24[19],_T_1003}; // @[Cat.scala 30:58]
  assign WallaceTree25_19_io_cin = WallaceTree25_18_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_20_io_n = {io_data_24[20],_T_1052}; // @[Cat.scala 30:58]
  assign WallaceTree25_20_io_cin = WallaceTree25_19_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_21_io_n = {io_data_24[21],_T_1101}; // @[Cat.scala 30:58]
  assign WallaceTree25_21_io_cin = WallaceTree25_20_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_22_io_n = {io_data_24[22],_T_1150}; // @[Cat.scala 30:58]
  assign WallaceTree25_22_io_cin = WallaceTree25_21_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_23_io_n = {io_data_24[23],_T_1199}; // @[Cat.scala 30:58]
  assign WallaceTree25_23_io_cin = WallaceTree25_22_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_24_io_n = {io_data_24[24],_T_1248}; // @[Cat.scala 30:58]
  assign WallaceTree25_24_io_cin = WallaceTree25_23_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_25_io_n = {io_data_24[25],_T_1297}; // @[Cat.scala 30:58]
  assign WallaceTree25_25_io_cin = WallaceTree25_24_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_26_io_n = {io_data_24[26],_T_1346}; // @[Cat.scala 30:58]
  assign WallaceTree25_26_io_cin = WallaceTree25_25_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_27_io_n = {io_data_24[27],_T_1395}; // @[Cat.scala 30:58]
  assign WallaceTree25_27_io_cin = WallaceTree25_26_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_28_io_n = {io_data_24[28],_T_1444}; // @[Cat.scala 30:58]
  assign WallaceTree25_28_io_cin = WallaceTree25_27_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_29_io_n = {io_data_24[29],_T_1493}; // @[Cat.scala 30:58]
  assign WallaceTree25_29_io_cin = WallaceTree25_28_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_30_io_n = {io_data_24[30],_T_1542}; // @[Cat.scala 30:58]
  assign WallaceTree25_30_io_cin = WallaceTree25_29_io_cout; // @[CNN_CONV.scala 161:{29,29}]
  assign WallaceTree25_31_io_n = {io_data_24[31],_T_1591}; // @[Cat.scala 30:58]
  assign WallaceTree25_31_io_cin = WallaceTree25_30_io_cout; // @[CNN_CONV.scala 161:{29,29}]
endmodule
module CNNConvSub25(
  input         clock,
  input         reset,
  input         io_conv_valid,
  input  [15:0] io_data_main_0,
  input  [15:0] io_data_main_1,
  input  [15:0] io_data_main_2,
  input  [15:0] io_data_main_3,
  input  [15:0] io_data_main_4,
  input  [15:0] io_data_main_5,
  input  [15:0] io_data_main_6,
  input  [15:0] io_data_main_7,
  input  [15:0] io_data_main_8,
  input  [15:0] io_data_main_9,
  input  [15:0] io_data_main_10,
  input  [15:0] io_data_main_11,
  input  [15:0] io_data_main_12,
  input  [15:0] io_data_main_13,
  input  [15:0] io_data_main_14,
  input  [15:0] io_data_main_15,
  input  [15:0] io_data_main_16,
  input  [15:0] io_data_main_17,
  input  [15:0] io_data_main_18,
  input  [15:0] io_data_main_19,
  input  [15:0] io_data_main_20,
  input  [15:0] io_data_main_21,
  input  [15:0] io_data_main_22,
  input  [15:0] io_data_main_23,
  input  [15:0] io_data_main_24,
  input  [7:0]  io_data_kernel_0,
  input  [7:0]  io_data_kernel_1,
  input  [7:0]  io_data_kernel_2,
  input  [7:0]  io_data_kernel_3,
  input  [7:0]  io_data_kernel_4,
  input  [7:0]  io_data_kernel_5,
  input  [7:0]  io_data_kernel_6,
  input  [7:0]  io_data_kernel_7,
  input  [7:0]  io_data_kernel_8,
  input  [7:0]  io_data_kernel_9,
  input  [7:0]  io_data_kernel_10,
  input  [7:0]  io_data_kernel_11,
  input  [7:0]  io_data_kernel_12,
  input  [7:0]  io_data_kernel_13,
  input  [7:0]  io_data_kernel_14,
  input  [7:0]  io_data_kernel_15,
  input  [7:0]  io_data_kernel_16,
  input  [7:0]  io_data_kernel_17,
  input  [7:0]  io_data_kernel_18,
  input  [7:0]  io_data_kernel_19,
  input  [7:0]  io_data_kernel_20,
  input  [7:0]  io_data_kernel_21,
  input  [7:0]  io_data_kernel_22,
  input  [7:0]  io_data_kernel_23,
  input  [7:0]  io_data_kernel_24,
  input  [3:0]  io_data_kernel_vwidth,
  output [31:0] io_data_res,
  output        io_data_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] BoothEncoderP_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_1_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_1_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_1_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_1_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_1_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_2_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_2_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_2_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_2_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_2_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_3_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_3_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_3_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_3_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_3_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_4_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_4_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_4_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_4_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_4_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_5_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_5_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_5_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_5_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_5_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_6_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_6_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_6_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_6_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_6_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_7_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_7_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_7_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_7_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_7_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_8_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_8_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_8_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_8_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_8_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_9_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_9_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_9_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_9_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_9_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_10_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_10_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_10_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_10_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_10_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_11_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_11_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_11_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_11_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_11_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_12_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_12_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_12_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_12_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_12_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_13_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_13_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_13_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_13_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_13_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_14_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_14_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_14_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_14_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_14_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_15_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_15_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_15_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_15_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_15_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_16_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_16_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_16_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_16_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_16_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_17_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_17_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_17_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_17_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_17_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_18_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_18_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_18_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_18_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_18_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_19_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_19_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_19_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_19_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_19_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_20_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_20_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_20_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_20_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_20_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_21_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_21_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_21_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_21_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_21_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_22_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_22_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_22_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_22_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_22_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_23_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_23_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_23_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_23_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_23_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_24_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_24_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_24_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_24_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_24_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_25_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_25_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_25_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_25_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_25_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_26_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_26_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_26_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_26_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_26_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_27_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_27_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_27_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_27_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_27_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_28_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_28_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_28_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_28_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_28_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_29_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_29_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_29_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_29_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_29_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_30_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_30_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_30_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_30_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_30_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_31_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_31_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_31_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_31_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_31_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_32_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_32_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_32_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_32_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_32_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_33_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_33_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_33_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_33_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_33_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_34_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_34_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_34_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_34_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_34_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_35_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_35_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_35_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_35_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_35_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_36_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_36_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_36_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_36_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_36_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_37_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_37_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_37_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_37_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_37_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_38_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_38_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_38_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_38_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_38_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_39_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_39_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_39_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_39_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_39_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_40_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_40_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_40_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_40_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_40_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_41_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_41_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_41_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_41_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_41_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_42_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_42_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_42_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_42_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_42_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_43_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_43_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_43_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_43_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_43_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_44_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_44_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_44_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_44_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_44_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_45_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_45_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_45_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_45_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_45_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_46_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_46_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_46_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_46_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_46_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_47_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_47_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_47_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_47_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_47_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_48_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_48_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_48_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_48_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_48_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_49_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_49_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_49_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_49_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_49_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_50_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_50_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_50_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_50_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_50_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_51_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_51_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_51_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_51_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_51_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_52_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_52_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_52_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_52_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_52_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_53_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_53_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_53_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_53_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_53_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_54_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_54_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_54_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_54_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_54_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_55_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_55_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_55_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_55_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_55_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_56_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_56_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_56_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_56_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_56_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_57_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_57_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_57_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_57_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_57_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_58_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_58_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_58_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_58_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_58_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_59_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_59_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_59_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_59_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_59_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_60_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_60_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_60_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_60_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_60_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_61_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_61_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_61_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_61_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_61_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_62_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_62_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_62_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_62_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_62_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_63_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_63_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_63_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_63_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_63_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_64_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_64_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_64_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_64_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_64_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_65_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_65_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_65_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_65_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_65_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_66_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_66_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_66_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_66_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_66_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_67_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_67_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_67_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_67_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_67_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_68_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_68_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_68_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_68_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_68_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_69_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_69_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_69_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_69_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_69_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_70_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_70_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_70_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_70_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_70_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_71_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_71_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_71_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_71_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_71_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_72_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_72_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_72_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_72_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_72_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_73_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_73_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_73_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_73_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_73_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_74_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_74_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_74_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_74_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_74_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_75_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_75_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_75_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_75_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_75_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_76_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_76_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_76_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_76_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_76_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_77_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_77_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_77_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_77_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_77_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_78_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_78_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_78_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_78_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_78_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_79_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_79_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_79_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_79_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_79_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_80_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_80_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_80_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_80_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_80_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_81_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_81_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_81_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_81_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_81_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_82_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_82_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_82_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_82_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_82_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_83_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_83_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_83_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_83_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_83_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_84_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_84_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_84_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_84_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_84_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_85_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_85_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_85_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_85_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_85_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_86_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_86_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_86_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_86_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_86_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_87_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_87_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_87_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_87_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_87_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_88_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_88_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_88_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_88_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_88_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_89_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_89_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_89_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_89_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_89_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_90_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_90_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_90_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_90_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_90_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_91_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_91_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_91_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_91_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_91_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_92_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_92_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_92_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_92_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_92_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_93_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_93_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_93_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_93_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_93_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_94_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_94_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_94_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_94_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_94_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_95_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_95_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_95_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_95_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_95_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_96_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_96_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_96_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_96_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_96_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_97_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_97_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_97_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_97_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_97_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_98_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_98_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_98_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_98_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_98_io_c; // @[CNN_CONV.scala 51:19]
  wire [2:0] BoothEncoderP_99_io_y; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_99_io_x; // @[CNN_CONV.scala 30:19]
  wire [31:0] BoothEncoderP_99_io_p; // @[CNN_CONV.scala 30:19]
  wire [2:0] BoothEncoderC_99_io_y; // @[CNN_CONV.scala 51:19]
  wire  BoothEncoderC_99_io_c; // @[CNN_CONV.scala 51:19]
  wire [31:0] WallaceAdder_io_data_0; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_1; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_2; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_3; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_4; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_5; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_6; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_7; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_8; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_9; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_10; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_11; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_12; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_13; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_14; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_15; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_16; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_17; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_18; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_19; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_20; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_21; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_22; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_23; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_data_24; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_0; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_1; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_2; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_3; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_4; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_5; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_6; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_7; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_8; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_9; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_10; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_11; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_12; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_13; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_14; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_15; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_16; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_17; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_18; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_19; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_20; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_21; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_22; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_23; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_io_cin_24; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_s; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_io_c; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_0; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_1; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_2; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_3; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_4; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_5; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_6; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_7; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_8; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_9; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_10; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_11; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_12; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_13; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_14; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_15; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_16; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_17; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_18; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_19; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_20; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_21; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_22; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_23; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_data_24; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_0; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_1; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_2; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_3; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_4; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_5; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_6; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_7; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_8; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_9; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_10; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_11; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_12; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_13; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_14; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_15; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_16; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_17; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_18; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_19; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_20; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_21; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_22; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_23; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_1_io_cin_24; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_s; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_1_io_c; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_0; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_1; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_2; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_3; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_4; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_5; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_6; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_7; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_8; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_9; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_10; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_11; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_12; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_13; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_14; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_15; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_16; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_17; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_18; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_19; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_20; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_21; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_22; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_23; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_data_24; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_0; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_1; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_2; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_3; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_4; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_5; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_6; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_7; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_8; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_9; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_10; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_11; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_12; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_13; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_14; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_15; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_16; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_17; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_18; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_19; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_20; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_21; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_22; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_23; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_2_io_cin_24; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_s; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_2_io_c; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_0; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_1; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_2; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_3; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_4; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_5; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_6; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_7; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_8; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_9; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_10; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_11; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_12; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_13; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_14; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_15; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_16; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_17; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_18; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_19; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_20; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_21; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_22; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_23; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_data_24; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_0; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_1; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_2; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_3; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_4; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_5; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_6; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_7; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_8; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_9; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_10; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_11; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_12; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_13; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_14; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_15; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_16; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_17; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_18; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_19; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_20; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_21; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_22; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_23; // @[CNN_CONV.scala 213:49]
  wire  WallaceAdder_3_io_cin_24; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_s; // @[CNN_CONV.scala 213:49]
  wire [31:0] WallaceAdder_3_io_c; // @[CNN_CONV.scala 213:49]
  wire [31:0] _T_2 = {16'h0,io_data_main_0}; // @[Cat.scala 30:58]
  wire [31:0] _T_7 = {16'h0,io_data_main_1}; // @[Cat.scala 30:58]
  wire [31:0] _T_12 = {16'h0,io_data_main_2}; // @[Cat.scala 30:58]
  wire [31:0] _T_17 = {16'h0,io_data_main_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_22 = {16'h0,io_data_main_4}; // @[Cat.scala 30:58]
  wire [31:0] _T_27 = {16'h0,io_data_main_5}; // @[Cat.scala 30:58]
  wire [31:0] _T_32 = {16'h0,io_data_main_6}; // @[Cat.scala 30:58]
  wire [31:0] _T_37 = {16'h0,io_data_main_7}; // @[Cat.scala 30:58]
  wire [31:0] _T_42 = {16'h0,io_data_main_8}; // @[Cat.scala 30:58]
  wire [31:0] _T_47 = {16'h0,io_data_main_9}; // @[Cat.scala 30:58]
  wire [31:0] _T_52 = {16'h0,io_data_main_10}; // @[Cat.scala 30:58]
  wire [31:0] _T_57 = {16'h0,io_data_main_11}; // @[Cat.scala 30:58]
  wire [31:0] _T_62 = {16'h0,io_data_main_12}; // @[Cat.scala 30:58]
  wire [31:0] _T_67 = {16'h0,io_data_main_13}; // @[Cat.scala 30:58]
  wire [31:0] _T_72 = {16'h0,io_data_main_14}; // @[Cat.scala 30:58]
  wire [31:0] _T_77 = {16'h0,io_data_main_15}; // @[Cat.scala 30:58]
  wire [31:0] _T_82 = {16'h0,io_data_main_16}; // @[Cat.scala 30:58]
  wire [31:0] _T_87 = {16'h0,io_data_main_17}; // @[Cat.scala 30:58]
  wire [31:0] _T_92 = {16'h0,io_data_main_18}; // @[Cat.scala 30:58]
  wire [31:0] _T_97 = {16'h0,io_data_main_19}; // @[Cat.scala 30:58]
  wire [31:0] _T_102 = {16'h0,io_data_main_20}; // @[Cat.scala 30:58]
  wire [31:0] _T_107 = {16'h0,io_data_main_21}; // @[Cat.scala 30:58]
  wire [31:0] _T_112 = {16'h0,io_data_main_22}; // @[Cat.scala 30:58]
  wire [31:0] _T_117 = {16'h0,io_data_main_23}; // @[Cat.scala 30:58]
  wire [31:0] _T_122 = {16'h0,io_data_main_24}; // @[Cat.scala 30:58]
  wire [33:0] _T_127 = {_T_2, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_131 = {_T_7, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_135 = {_T_12, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_139 = {_T_17, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_143 = {_T_22, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_147 = {_T_27, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_151 = {_T_32, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_155 = {_T_37, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_159 = {_T_42, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_163 = {_T_47, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_167 = {_T_52, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_171 = {_T_57, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_175 = {_T_62, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_179 = {_T_67, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_183 = {_T_72, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_187 = {_T_77, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_191 = {_T_82, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_195 = {_T_87, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_199 = {_T_92, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_203 = {_T_97, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_207 = {_T_102, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_211 = {_T_107, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_215 = {_T_112, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_219 = {_T_117, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [33:0] _T_223 = {_T_122, 2'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_227 = {_T_2, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_231 = {_T_7, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_235 = {_T_12, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_239 = {_T_17, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_243 = {_T_22, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_247 = {_T_27, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_251 = {_T_32, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_255 = {_T_37, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_259 = {_T_42, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_263 = {_T_47, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_267 = {_T_52, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_271 = {_T_57, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_275 = {_T_62, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_279 = {_T_67, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_283 = {_T_72, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_287 = {_T_77, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_291 = {_T_82, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_295 = {_T_87, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_299 = {_T_92, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_303 = {_T_97, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_307 = {_T_102, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_311 = {_T_107, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_315 = {_T_112, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_319 = {_T_117, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [35:0] _T_323 = {_T_122, 4'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_327 = {_T_2, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_331 = {_T_7, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_335 = {_T_12, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_339 = {_T_17, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_343 = {_T_22, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_347 = {_T_27, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_351 = {_T_32, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_355 = {_T_37, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_359 = {_T_42, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_363 = {_T_47, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_367 = {_T_52, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_371 = {_T_57, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_375 = {_T_62, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_379 = {_T_67, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_383 = {_T_72, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_387 = {_T_77, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_391 = {_T_82, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_395 = {_T_87, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_399 = {_T_92, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_403 = {_T_97, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_407 = {_T_102, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_411 = {_T_107, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_415 = {_T_112, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_419 = {_T_117, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [37:0] _T_423 = {_T_122, 6'h0}; // @[CNN_CONV.scala 206:103]
  wire [31:0] wallace_adder_0_s = WallaceAdder_io_s; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] wallace_adder_0_c = WallaceAdder_io_c; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] res_int21 = wallace_adder_0_s + wallace_adder_0_c; // @[CNN_CONV.scala 223:28]
  reg  state; // @[CNN_CONV.scala 228:22]
  wire  _T_426 = ~state; // @[CNN_CONV.scala 229:46]
  wire  stage2_valid = io_conv_valid & ~state & (io_data_kernel_vwidth[3] | io_data_kernel_vwidth[2]); // @[CNN_CONV.scala 229:60]
  wire  _GEN_0 = stage2_valid | state; // @[CNN_CONV.scala 228:22 232:{29,37}]
  reg [31:0] out_s_reg_0; // @[CNN_CONV.scala 238:26]
  reg [31:0] out_s_reg_1; // @[CNN_CONV.scala 238:26]
  reg [31:0] out_s_reg_2; // @[CNN_CONV.scala 238:26]
  reg [31:0] out_s_reg_3; // @[CNN_CONV.scala 238:26]
  reg [31:0] out_c_reg_0; // @[CNN_CONV.scala 239:26]
  reg [31:0] out_c_reg_1; // @[CNN_CONV.scala 239:26]
  reg [31:0] out_c_reg_2; // @[CNN_CONV.scala 239:26]
  reg [31:0] out_c_reg_3; // @[CNN_CONV.scala 239:26]
  wire [31:0] wallace_adder_1_s = WallaceAdder_1_io_s; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] wallace_adder_2_s = WallaceAdder_2_io_s; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] wallace_adder_3_s = WallaceAdder_3_io_s; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] wallace_adder_1_c = WallaceAdder_1_io_c; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] wallace_adder_2_c = WallaceAdder_2_io_c; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] wallace_adder_3_c = WallaceAdder_3_io_c; // @[CNN_CONV.scala 213:{30,30}]
  wire [31:0] _T_434 = out_s_reg_0 + out_s_reg_1; // @[CNN_CONV.scala 243:37]
  wire [31:0] _T_436 = _T_434 + out_s_reg_2; // @[CNN_CONV.scala 243:37]
  wire [31:0] _T_438 = _T_436 + out_s_reg_3; // @[CNN_CONV.scala 243:37]
  wire [31:0] _T_440 = out_c_reg_0 + out_c_reg_1; // @[CNN_CONV.scala 243:63]
  wire [31:0] _T_442 = _T_440 + out_c_reg_2; // @[CNN_CONV.scala 243:63]
  wire [31:0] _T_444 = _T_442 + out_c_reg_3; // @[CNN_CONV.scala 243:63]
  wire [31:0] res_int8 = _T_438 + _T_444; // @[CNN_CONV.scala 243:42]
  wire [31:0] _T_449 = _T_434 + out_c_reg_0; // @[CNN_CONV.scala 244:46]
  wire [31:0] res_int4 = _T_449 + out_c_reg_1; // @[CNN_CONV.scala 244:61]
  wire [31:0] _T_453 = io_data_kernel_vwidth[3] ? res_int8 : res_int4; // @[CNN_CONV.scala 247:46]
  BoothEncoderP BoothEncoderP ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_io_y),
    .io_x(BoothEncoderP_io_x),
    .io_p(BoothEncoderP_io_p)
  );
  BoothEncoderC BoothEncoderC ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_io_y),
    .io_c(BoothEncoderC_io_c)
  );
  BoothEncoderP BoothEncoderP_1 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_1_io_y),
    .io_x(BoothEncoderP_1_io_x),
    .io_p(BoothEncoderP_1_io_p)
  );
  BoothEncoderC BoothEncoderC_1 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_1_io_y),
    .io_c(BoothEncoderC_1_io_c)
  );
  BoothEncoderP BoothEncoderP_2 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_2_io_y),
    .io_x(BoothEncoderP_2_io_x),
    .io_p(BoothEncoderP_2_io_p)
  );
  BoothEncoderC BoothEncoderC_2 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_2_io_y),
    .io_c(BoothEncoderC_2_io_c)
  );
  BoothEncoderP BoothEncoderP_3 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_3_io_y),
    .io_x(BoothEncoderP_3_io_x),
    .io_p(BoothEncoderP_3_io_p)
  );
  BoothEncoderC BoothEncoderC_3 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_3_io_y),
    .io_c(BoothEncoderC_3_io_c)
  );
  BoothEncoderP BoothEncoderP_4 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_4_io_y),
    .io_x(BoothEncoderP_4_io_x),
    .io_p(BoothEncoderP_4_io_p)
  );
  BoothEncoderC BoothEncoderC_4 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_4_io_y),
    .io_c(BoothEncoderC_4_io_c)
  );
  BoothEncoderP BoothEncoderP_5 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_5_io_y),
    .io_x(BoothEncoderP_5_io_x),
    .io_p(BoothEncoderP_5_io_p)
  );
  BoothEncoderC BoothEncoderC_5 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_5_io_y),
    .io_c(BoothEncoderC_5_io_c)
  );
  BoothEncoderP BoothEncoderP_6 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_6_io_y),
    .io_x(BoothEncoderP_6_io_x),
    .io_p(BoothEncoderP_6_io_p)
  );
  BoothEncoderC BoothEncoderC_6 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_6_io_y),
    .io_c(BoothEncoderC_6_io_c)
  );
  BoothEncoderP BoothEncoderP_7 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_7_io_y),
    .io_x(BoothEncoderP_7_io_x),
    .io_p(BoothEncoderP_7_io_p)
  );
  BoothEncoderC BoothEncoderC_7 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_7_io_y),
    .io_c(BoothEncoderC_7_io_c)
  );
  BoothEncoderP BoothEncoderP_8 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_8_io_y),
    .io_x(BoothEncoderP_8_io_x),
    .io_p(BoothEncoderP_8_io_p)
  );
  BoothEncoderC BoothEncoderC_8 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_8_io_y),
    .io_c(BoothEncoderC_8_io_c)
  );
  BoothEncoderP BoothEncoderP_9 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_9_io_y),
    .io_x(BoothEncoderP_9_io_x),
    .io_p(BoothEncoderP_9_io_p)
  );
  BoothEncoderC BoothEncoderC_9 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_9_io_y),
    .io_c(BoothEncoderC_9_io_c)
  );
  BoothEncoderP BoothEncoderP_10 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_10_io_y),
    .io_x(BoothEncoderP_10_io_x),
    .io_p(BoothEncoderP_10_io_p)
  );
  BoothEncoderC BoothEncoderC_10 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_10_io_y),
    .io_c(BoothEncoderC_10_io_c)
  );
  BoothEncoderP BoothEncoderP_11 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_11_io_y),
    .io_x(BoothEncoderP_11_io_x),
    .io_p(BoothEncoderP_11_io_p)
  );
  BoothEncoderC BoothEncoderC_11 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_11_io_y),
    .io_c(BoothEncoderC_11_io_c)
  );
  BoothEncoderP BoothEncoderP_12 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_12_io_y),
    .io_x(BoothEncoderP_12_io_x),
    .io_p(BoothEncoderP_12_io_p)
  );
  BoothEncoderC BoothEncoderC_12 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_12_io_y),
    .io_c(BoothEncoderC_12_io_c)
  );
  BoothEncoderP BoothEncoderP_13 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_13_io_y),
    .io_x(BoothEncoderP_13_io_x),
    .io_p(BoothEncoderP_13_io_p)
  );
  BoothEncoderC BoothEncoderC_13 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_13_io_y),
    .io_c(BoothEncoderC_13_io_c)
  );
  BoothEncoderP BoothEncoderP_14 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_14_io_y),
    .io_x(BoothEncoderP_14_io_x),
    .io_p(BoothEncoderP_14_io_p)
  );
  BoothEncoderC BoothEncoderC_14 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_14_io_y),
    .io_c(BoothEncoderC_14_io_c)
  );
  BoothEncoderP BoothEncoderP_15 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_15_io_y),
    .io_x(BoothEncoderP_15_io_x),
    .io_p(BoothEncoderP_15_io_p)
  );
  BoothEncoderC BoothEncoderC_15 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_15_io_y),
    .io_c(BoothEncoderC_15_io_c)
  );
  BoothEncoderP BoothEncoderP_16 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_16_io_y),
    .io_x(BoothEncoderP_16_io_x),
    .io_p(BoothEncoderP_16_io_p)
  );
  BoothEncoderC BoothEncoderC_16 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_16_io_y),
    .io_c(BoothEncoderC_16_io_c)
  );
  BoothEncoderP BoothEncoderP_17 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_17_io_y),
    .io_x(BoothEncoderP_17_io_x),
    .io_p(BoothEncoderP_17_io_p)
  );
  BoothEncoderC BoothEncoderC_17 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_17_io_y),
    .io_c(BoothEncoderC_17_io_c)
  );
  BoothEncoderP BoothEncoderP_18 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_18_io_y),
    .io_x(BoothEncoderP_18_io_x),
    .io_p(BoothEncoderP_18_io_p)
  );
  BoothEncoderC BoothEncoderC_18 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_18_io_y),
    .io_c(BoothEncoderC_18_io_c)
  );
  BoothEncoderP BoothEncoderP_19 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_19_io_y),
    .io_x(BoothEncoderP_19_io_x),
    .io_p(BoothEncoderP_19_io_p)
  );
  BoothEncoderC BoothEncoderC_19 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_19_io_y),
    .io_c(BoothEncoderC_19_io_c)
  );
  BoothEncoderP BoothEncoderP_20 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_20_io_y),
    .io_x(BoothEncoderP_20_io_x),
    .io_p(BoothEncoderP_20_io_p)
  );
  BoothEncoderC BoothEncoderC_20 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_20_io_y),
    .io_c(BoothEncoderC_20_io_c)
  );
  BoothEncoderP BoothEncoderP_21 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_21_io_y),
    .io_x(BoothEncoderP_21_io_x),
    .io_p(BoothEncoderP_21_io_p)
  );
  BoothEncoderC BoothEncoderC_21 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_21_io_y),
    .io_c(BoothEncoderC_21_io_c)
  );
  BoothEncoderP BoothEncoderP_22 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_22_io_y),
    .io_x(BoothEncoderP_22_io_x),
    .io_p(BoothEncoderP_22_io_p)
  );
  BoothEncoderC BoothEncoderC_22 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_22_io_y),
    .io_c(BoothEncoderC_22_io_c)
  );
  BoothEncoderP BoothEncoderP_23 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_23_io_y),
    .io_x(BoothEncoderP_23_io_x),
    .io_p(BoothEncoderP_23_io_p)
  );
  BoothEncoderC BoothEncoderC_23 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_23_io_y),
    .io_c(BoothEncoderC_23_io_c)
  );
  BoothEncoderP BoothEncoderP_24 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_24_io_y),
    .io_x(BoothEncoderP_24_io_x),
    .io_p(BoothEncoderP_24_io_p)
  );
  BoothEncoderC BoothEncoderC_24 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_24_io_y),
    .io_c(BoothEncoderC_24_io_c)
  );
  BoothEncoderP BoothEncoderP_25 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_25_io_y),
    .io_x(BoothEncoderP_25_io_x),
    .io_p(BoothEncoderP_25_io_p)
  );
  BoothEncoderC BoothEncoderC_25 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_25_io_y),
    .io_c(BoothEncoderC_25_io_c)
  );
  BoothEncoderP BoothEncoderP_26 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_26_io_y),
    .io_x(BoothEncoderP_26_io_x),
    .io_p(BoothEncoderP_26_io_p)
  );
  BoothEncoderC BoothEncoderC_26 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_26_io_y),
    .io_c(BoothEncoderC_26_io_c)
  );
  BoothEncoderP BoothEncoderP_27 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_27_io_y),
    .io_x(BoothEncoderP_27_io_x),
    .io_p(BoothEncoderP_27_io_p)
  );
  BoothEncoderC BoothEncoderC_27 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_27_io_y),
    .io_c(BoothEncoderC_27_io_c)
  );
  BoothEncoderP BoothEncoderP_28 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_28_io_y),
    .io_x(BoothEncoderP_28_io_x),
    .io_p(BoothEncoderP_28_io_p)
  );
  BoothEncoderC BoothEncoderC_28 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_28_io_y),
    .io_c(BoothEncoderC_28_io_c)
  );
  BoothEncoderP BoothEncoderP_29 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_29_io_y),
    .io_x(BoothEncoderP_29_io_x),
    .io_p(BoothEncoderP_29_io_p)
  );
  BoothEncoderC BoothEncoderC_29 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_29_io_y),
    .io_c(BoothEncoderC_29_io_c)
  );
  BoothEncoderP BoothEncoderP_30 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_30_io_y),
    .io_x(BoothEncoderP_30_io_x),
    .io_p(BoothEncoderP_30_io_p)
  );
  BoothEncoderC BoothEncoderC_30 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_30_io_y),
    .io_c(BoothEncoderC_30_io_c)
  );
  BoothEncoderP BoothEncoderP_31 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_31_io_y),
    .io_x(BoothEncoderP_31_io_x),
    .io_p(BoothEncoderP_31_io_p)
  );
  BoothEncoderC BoothEncoderC_31 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_31_io_y),
    .io_c(BoothEncoderC_31_io_c)
  );
  BoothEncoderP BoothEncoderP_32 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_32_io_y),
    .io_x(BoothEncoderP_32_io_x),
    .io_p(BoothEncoderP_32_io_p)
  );
  BoothEncoderC BoothEncoderC_32 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_32_io_y),
    .io_c(BoothEncoderC_32_io_c)
  );
  BoothEncoderP BoothEncoderP_33 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_33_io_y),
    .io_x(BoothEncoderP_33_io_x),
    .io_p(BoothEncoderP_33_io_p)
  );
  BoothEncoderC BoothEncoderC_33 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_33_io_y),
    .io_c(BoothEncoderC_33_io_c)
  );
  BoothEncoderP BoothEncoderP_34 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_34_io_y),
    .io_x(BoothEncoderP_34_io_x),
    .io_p(BoothEncoderP_34_io_p)
  );
  BoothEncoderC BoothEncoderC_34 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_34_io_y),
    .io_c(BoothEncoderC_34_io_c)
  );
  BoothEncoderP BoothEncoderP_35 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_35_io_y),
    .io_x(BoothEncoderP_35_io_x),
    .io_p(BoothEncoderP_35_io_p)
  );
  BoothEncoderC BoothEncoderC_35 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_35_io_y),
    .io_c(BoothEncoderC_35_io_c)
  );
  BoothEncoderP BoothEncoderP_36 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_36_io_y),
    .io_x(BoothEncoderP_36_io_x),
    .io_p(BoothEncoderP_36_io_p)
  );
  BoothEncoderC BoothEncoderC_36 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_36_io_y),
    .io_c(BoothEncoderC_36_io_c)
  );
  BoothEncoderP BoothEncoderP_37 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_37_io_y),
    .io_x(BoothEncoderP_37_io_x),
    .io_p(BoothEncoderP_37_io_p)
  );
  BoothEncoderC BoothEncoderC_37 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_37_io_y),
    .io_c(BoothEncoderC_37_io_c)
  );
  BoothEncoderP BoothEncoderP_38 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_38_io_y),
    .io_x(BoothEncoderP_38_io_x),
    .io_p(BoothEncoderP_38_io_p)
  );
  BoothEncoderC BoothEncoderC_38 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_38_io_y),
    .io_c(BoothEncoderC_38_io_c)
  );
  BoothEncoderP BoothEncoderP_39 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_39_io_y),
    .io_x(BoothEncoderP_39_io_x),
    .io_p(BoothEncoderP_39_io_p)
  );
  BoothEncoderC BoothEncoderC_39 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_39_io_y),
    .io_c(BoothEncoderC_39_io_c)
  );
  BoothEncoderP BoothEncoderP_40 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_40_io_y),
    .io_x(BoothEncoderP_40_io_x),
    .io_p(BoothEncoderP_40_io_p)
  );
  BoothEncoderC BoothEncoderC_40 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_40_io_y),
    .io_c(BoothEncoderC_40_io_c)
  );
  BoothEncoderP BoothEncoderP_41 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_41_io_y),
    .io_x(BoothEncoderP_41_io_x),
    .io_p(BoothEncoderP_41_io_p)
  );
  BoothEncoderC BoothEncoderC_41 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_41_io_y),
    .io_c(BoothEncoderC_41_io_c)
  );
  BoothEncoderP BoothEncoderP_42 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_42_io_y),
    .io_x(BoothEncoderP_42_io_x),
    .io_p(BoothEncoderP_42_io_p)
  );
  BoothEncoderC BoothEncoderC_42 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_42_io_y),
    .io_c(BoothEncoderC_42_io_c)
  );
  BoothEncoderP BoothEncoderP_43 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_43_io_y),
    .io_x(BoothEncoderP_43_io_x),
    .io_p(BoothEncoderP_43_io_p)
  );
  BoothEncoderC BoothEncoderC_43 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_43_io_y),
    .io_c(BoothEncoderC_43_io_c)
  );
  BoothEncoderP BoothEncoderP_44 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_44_io_y),
    .io_x(BoothEncoderP_44_io_x),
    .io_p(BoothEncoderP_44_io_p)
  );
  BoothEncoderC BoothEncoderC_44 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_44_io_y),
    .io_c(BoothEncoderC_44_io_c)
  );
  BoothEncoderP BoothEncoderP_45 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_45_io_y),
    .io_x(BoothEncoderP_45_io_x),
    .io_p(BoothEncoderP_45_io_p)
  );
  BoothEncoderC BoothEncoderC_45 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_45_io_y),
    .io_c(BoothEncoderC_45_io_c)
  );
  BoothEncoderP BoothEncoderP_46 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_46_io_y),
    .io_x(BoothEncoderP_46_io_x),
    .io_p(BoothEncoderP_46_io_p)
  );
  BoothEncoderC BoothEncoderC_46 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_46_io_y),
    .io_c(BoothEncoderC_46_io_c)
  );
  BoothEncoderP BoothEncoderP_47 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_47_io_y),
    .io_x(BoothEncoderP_47_io_x),
    .io_p(BoothEncoderP_47_io_p)
  );
  BoothEncoderC BoothEncoderC_47 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_47_io_y),
    .io_c(BoothEncoderC_47_io_c)
  );
  BoothEncoderP BoothEncoderP_48 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_48_io_y),
    .io_x(BoothEncoderP_48_io_x),
    .io_p(BoothEncoderP_48_io_p)
  );
  BoothEncoderC BoothEncoderC_48 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_48_io_y),
    .io_c(BoothEncoderC_48_io_c)
  );
  BoothEncoderP BoothEncoderP_49 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_49_io_y),
    .io_x(BoothEncoderP_49_io_x),
    .io_p(BoothEncoderP_49_io_p)
  );
  BoothEncoderC BoothEncoderC_49 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_49_io_y),
    .io_c(BoothEncoderC_49_io_c)
  );
  BoothEncoderP BoothEncoderP_50 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_50_io_y),
    .io_x(BoothEncoderP_50_io_x),
    .io_p(BoothEncoderP_50_io_p)
  );
  BoothEncoderC BoothEncoderC_50 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_50_io_y),
    .io_c(BoothEncoderC_50_io_c)
  );
  BoothEncoderP BoothEncoderP_51 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_51_io_y),
    .io_x(BoothEncoderP_51_io_x),
    .io_p(BoothEncoderP_51_io_p)
  );
  BoothEncoderC BoothEncoderC_51 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_51_io_y),
    .io_c(BoothEncoderC_51_io_c)
  );
  BoothEncoderP BoothEncoderP_52 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_52_io_y),
    .io_x(BoothEncoderP_52_io_x),
    .io_p(BoothEncoderP_52_io_p)
  );
  BoothEncoderC BoothEncoderC_52 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_52_io_y),
    .io_c(BoothEncoderC_52_io_c)
  );
  BoothEncoderP BoothEncoderP_53 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_53_io_y),
    .io_x(BoothEncoderP_53_io_x),
    .io_p(BoothEncoderP_53_io_p)
  );
  BoothEncoderC BoothEncoderC_53 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_53_io_y),
    .io_c(BoothEncoderC_53_io_c)
  );
  BoothEncoderP BoothEncoderP_54 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_54_io_y),
    .io_x(BoothEncoderP_54_io_x),
    .io_p(BoothEncoderP_54_io_p)
  );
  BoothEncoderC BoothEncoderC_54 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_54_io_y),
    .io_c(BoothEncoderC_54_io_c)
  );
  BoothEncoderP BoothEncoderP_55 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_55_io_y),
    .io_x(BoothEncoderP_55_io_x),
    .io_p(BoothEncoderP_55_io_p)
  );
  BoothEncoderC BoothEncoderC_55 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_55_io_y),
    .io_c(BoothEncoderC_55_io_c)
  );
  BoothEncoderP BoothEncoderP_56 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_56_io_y),
    .io_x(BoothEncoderP_56_io_x),
    .io_p(BoothEncoderP_56_io_p)
  );
  BoothEncoderC BoothEncoderC_56 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_56_io_y),
    .io_c(BoothEncoderC_56_io_c)
  );
  BoothEncoderP BoothEncoderP_57 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_57_io_y),
    .io_x(BoothEncoderP_57_io_x),
    .io_p(BoothEncoderP_57_io_p)
  );
  BoothEncoderC BoothEncoderC_57 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_57_io_y),
    .io_c(BoothEncoderC_57_io_c)
  );
  BoothEncoderP BoothEncoderP_58 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_58_io_y),
    .io_x(BoothEncoderP_58_io_x),
    .io_p(BoothEncoderP_58_io_p)
  );
  BoothEncoderC BoothEncoderC_58 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_58_io_y),
    .io_c(BoothEncoderC_58_io_c)
  );
  BoothEncoderP BoothEncoderP_59 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_59_io_y),
    .io_x(BoothEncoderP_59_io_x),
    .io_p(BoothEncoderP_59_io_p)
  );
  BoothEncoderC BoothEncoderC_59 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_59_io_y),
    .io_c(BoothEncoderC_59_io_c)
  );
  BoothEncoderP BoothEncoderP_60 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_60_io_y),
    .io_x(BoothEncoderP_60_io_x),
    .io_p(BoothEncoderP_60_io_p)
  );
  BoothEncoderC BoothEncoderC_60 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_60_io_y),
    .io_c(BoothEncoderC_60_io_c)
  );
  BoothEncoderP BoothEncoderP_61 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_61_io_y),
    .io_x(BoothEncoderP_61_io_x),
    .io_p(BoothEncoderP_61_io_p)
  );
  BoothEncoderC BoothEncoderC_61 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_61_io_y),
    .io_c(BoothEncoderC_61_io_c)
  );
  BoothEncoderP BoothEncoderP_62 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_62_io_y),
    .io_x(BoothEncoderP_62_io_x),
    .io_p(BoothEncoderP_62_io_p)
  );
  BoothEncoderC BoothEncoderC_62 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_62_io_y),
    .io_c(BoothEncoderC_62_io_c)
  );
  BoothEncoderP BoothEncoderP_63 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_63_io_y),
    .io_x(BoothEncoderP_63_io_x),
    .io_p(BoothEncoderP_63_io_p)
  );
  BoothEncoderC BoothEncoderC_63 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_63_io_y),
    .io_c(BoothEncoderC_63_io_c)
  );
  BoothEncoderP BoothEncoderP_64 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_64_io_y),
    .io_x(BoothEncoderP_64_io_x),
    .io_p(BoothEncoderP_64_io_p)
  );
  BoothEncoderC BoothEncoderC_64 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_64_io_y),
    .io_c(BoothEncoderC_64_io_c)
  );
  BoothEncoderP BoothEncoderP_65 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_65_io_y),
    .io_x(BoothEncoderP_65_io_x),
    .io_p(BoothEncoderP_65_io_p)
  );
  BoothEncoderC BoothEncoderC_65 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_65_io_y),
    .io_c(BoothEncoderC_65_io_c)
  );
  BoothEncoderP BoothEncoderP_66 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_66_io_y),
    .io_x(BoothEncoderP_66_io_x),
    .io_p(BoothEncoderP_66_io_p)
  );
  BoothEncoderC BoothEncoderC_66 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_66_io_y),
    .io_c(BoothEncoderC_66_io_c)
  );
  BoothEncoderP BoothEncoderP_67 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_67_io_y),
    .io_x(BoothEncoderP_67_io_x),
    .io_p(BoothEncoderP_67_io_p)
  );
  BoothEncoderC BoothEncoderC_67 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_67_io_y),
    .io_c(BoothEncoderC_67_io_c)
  );
  BoothEncoderP BoothEncoderP_68 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_68_io_y),
    .io_x(BoothEncoderP_68_io_x),
    .io_p(BoothEncoderP_68_io_p)
  );
  BoothEncoderC BoothEncoderC_68 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_68_io_y),
    .io_c(BoothEncoderC_68_io_c)
  );
  BoothEncoderP BoothEncoderP_69 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_69_io_y),
    .io_x(BoothEncoderP_69_io_x),
    .io_p(BoothEncoderP_69_io_p)
  );
  BoothEncoderC BoothEncoderC_69 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_69_io_y),
    .io_c(BoothEncoderC_69_io_c)
  );
  BoothEncoderP BoothEncoderP_70 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_70_io_y),
    .io_x(BoothEncoderP_70_io_x),
    .io_p(BoothEncoderP_70_io_p)
  );
  BoothEncoderC BoothEncoderC_70 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_70_io_y),
    .io_c(BoothEncoderC_70_io_c)
  );
  BoothEncoderP BoothEncoderP_71 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_71_io_y),
    .io_x(BoothEncoderP_71_io_x),
    .io_p(BoothEncoderP_71_io_p)
  );
  BoothEncoderC BoothEncoderC_71 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_71_io_y),
    .io_c(BoothEncoderC_71_io_c)
  );
  BoothEncoderP BoothEncoderP_72 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_72_io_y),
    .io_x(BoothEncoderP_72_io_x),
    .io_p(BoothEncoderP_72_io_p)
  );
  BoothEncoderC BoothEncoderC_72 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_72_io_y),
    .io_c(BoothEncoderC_72_io_c)
  );
  BoothEncoderP BoothEncoderP_73 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_73_io_y),
    .io_x(BoothEncoderP_73_io_x),
    .io_p(BoothEncoderP_73_io_p)
  );
  BoothEncoderC BoothEncoderC_73 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_73_io_y),
    .io_c(BoothEncoderC_73_io_c)
  );
  BoothEncoderP BoothEncoderP_74 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_74_io_y),
    .io_x(BoothEncoderP_74_io_x),
    .io_p(BoothEncoderP_74_io_p)
  );
  BoothEncoderC BoothEncoderC_74 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_74_io_y),
    .io_c(BoothEncoderC_74_io_c)
  );
  BoothEncoderP BoothEncoderP_75 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_75_io_y),
    .io_x(BoothEncoderP_75_io_x),
    .io_p(BoothEncoderP_75_io_p)
  );
  BoothEncoderC BoothEncoderC_75 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_75_io_y),
    .io_c(BoothEncoderC_75_io_c)
  );
  BoothEncoderP BoothEncoderP_76 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_76_io_y),
    .io_x(BoothEncoderP_76_io_x),
    .io_p(BoothEncoderP_76_io_p)
  );
  BoothEncoderC BoothEncoderC_76 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_76_io_y),
    .io_c(BoothEncoderC_76_io_c)
  );
  BoothEncoderP BoothEncoderP_77 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_77_io_y),
    .io_x(BoothEncoderP_77_io_x),
    .io_p(BoothEncoderP_77_io_p)
  );
  BoothEncoderC BoothEncoderC_77 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_77_io_y),
    .io_c(BoothEncoderC_77_io_c)
  );
  BoothEncoderP BoothEncoderP_78 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_78_io_y),
    .io_x(BoothEncoderP_78_io_x),
    .io_p(BoothEncoderP_78_io_p)
  );
  BoothEncoderC BoothEncoderC_78 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_78_io_y),
    .io_c(BoothEncoderC_78_io_c)
  );
  BoothEncoderP BoothEncoderP_79 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_79_io_y),
    .io_x(BoothEncoderP_79_io_x),
    .io_p(BoothEncoderP_79_io_p)
  );
  BoothEncoderC BoothEncoderC_79 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_79_io_y),
    .io_c(BoothEncoderC_79_io_c)
  );
  BoothEncoderP BoothEncoderP_80 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_80_io_y),
    .io_x(BoothEncoderP_80_io_x),
    .io_p(BoothEncoderP_80_io_p)
  );
  BoothEncoderC BoothEncoderC_80 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_80_io_y),
    .io_c(BoothEncoderC_80_io_c)
  );
  BoothEncoderP BoothEncoderP_81 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_81_io_y),
    .io_x(BoothEncoderP_81_io_x),
    .io_p(BoothEncoderP_81_io_p)
  );
  BoothEncoderC BoothEncoderC_81 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_81_io_y),
    .io_c(BoothEncoderC_81_io_c)
  );
  BoothEncoderP BoothEncoderP_82 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_82_io_y),
    .io_x(BoothEncoderP_82_io_x),
    .io_p(BoothEncoderP_82_io_p)
  );
  BoothEncoderC BoothEncoderC_82 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_82_io_y),
    .io_c(BoothEncoderC_82_io_c)
  );
  BoothEncoderP BoothEncoderP_83 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_83_io_y),
    .io_x(BoothEncoderP_83_io_x),
    .io_p(BoothEncoderP_83_io_p)
  );
  BoothEncoderC BoothEncoderC_83 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_83_io_y),
    .io_c(BoothEncoderC_83_io_c)
  );
  BoothEncoderP BoothEncoderP_84 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_84_io_y),
    .io_x(BoothEncoderP_84_io_x),
    .io_p(BoothEncoderP_84_io_p)
  );
  BoothEncoderC BoothEncoderC_84 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_84_io_y),
    .io_c(BoothEncoderC_84_io_c)
  );
  BoothEncoderP BoothEncoderP_85 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_85_io_y),
    .io_x(BoothEncoderP_85_io_x),
    .io_p(BoothEncoderP_85_io_p)
  );
  BoothEncoderC BoothEncoderC_85 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_85_io_y),
    .io_c(BoothEncoderC_85_io_c)
  );
  BoothEncoderP BoothEncoderP_86 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_86_io_y),
    .io_x(BoothEncoderP_86_io_x),
    .io_p(BoothEncoderP_86_io_p)
  );
  BoothEncoderC BoothEncoderC_86 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_86_io_y),
    .io_c(BoothEncoderC_86_io_c)
  );
  BoothEncoderP BoothEncoderP_87 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_87_io_y),
    .io_x(BoothEncoderP_87_io_x),
    .io_p(BoothEncoderP_87_io_p)
  );
  BoothEncoderC BoothEncoderC_87 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_87_io_y),
    .io_c(BoothEncoderC_87_io_c)
  );
  BoothEncoderP BoothEncoderP_88 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_88_io_y),
    .io_x(BoothEncoderP_88_io_x),
    .io_p(BoothEncoderP_88_io_p)
  );
  BoothEncoderC BoothEncoderC_88 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_88_io_y),
    .io_c(BoothEncoderC_88_io_c)
  );
  BoothEncoderP BoothEncoderP_89 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_89_io_y),
    .io_x(BoothEncoderP_89_io_x),
    .io_p(BoothEncoderP_89_io_p)
  );
  BoothEncoderC BoothEncoderC_89 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_89_io_y),
    .io_c(BoothEncoderC_89_io_c)
  );
  BoothEncoderP BoothEncoderP_90 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_90_io_y),
    .io_x(BoothEncoderP_90_io_x),
    .io_p(BoothEncoderP_90_io_p)
  );
  BoothEncoderC BoothEncoderC_90 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_90_io_y),
    .io_c(BoothEncoderC_90_io_c)
  );
  BoothEncoderP BoothEncoderP_91 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_91_io_y),
    .io_x(BoothEncoderP_91_io_x),
    .io_p(BoothEncoderP_91_io_p)
  );
  BoothEncoderC BoothEncoderC_91 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_91_io_y),
    .io_c(BoothEncoderC_91_io_c)
  );
  BoothEncoderP BoothEncoderP_92 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_92_io_y),
    .io_x(BoothEncoderP_92_io_x),
    .io_p(BoothEncoderP_92_io_p)
  );
  BoothEncoderC BoothEncoderC_92 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_92_io_y),
    .io_c(BoothEncoderC_92_io_c)
  );
  BoothEncoderP BoothEncoderP_93 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_93_io_y),
    .io_x(BoothEncoderP_93_io_x),
    .io_p(BoothEncoderP_93_io_p)
  );
  BoothEncoderC BoothEncoderC_93 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_93_io_y),
    .io_c(BoothEncoderC_93_io_c)
  );
  BoothEncoderP BoothEncoderP_94 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_94_io_y),
    .io_x(BoothEncoderP_94_io_x),
    .io_p(BoothEncoderP_94_io_p)
  );
  BoothEncoderC BoothEncoderC_94 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_94_io_y),
    .io_c(BoothEncoderC_94_io_c)
  );
  BoothEncoderP BoothEncoderP_95 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_95_io_y),
    .io_x(BoothEncoderP_95_io_x),
    .io_p(BoothEncoderP_95_io_p)
  );
  BoothEncoderC BoothEncoderC_95 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_95_io_y),
    .io_c(BoothEncoderC_95_io_c)
  );
  BoothEncoderP BoothEncoderP_96 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_96_io_y),
    .io_x(BoothEncoderP_96_io_x),
    .io_p(BoothEncoderP_96_io_p)
  );
  BoothEncoderC BoothEncoderC_96 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_96_io_y),
    .io_c(BoothEncoderC_96_io_c)
  );
  BoothEncoderP BoothEncoderP_97 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_97_io_y),
    .io_x(BoothEncoderP_97_io_x),
    .io_p(BoothEncoderP_97_io_p)
  );
  BoothEncoderC BoothEncoderC_97 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_97_io_y),
    .io_c(BoothEncoderC_97_io_c)
  );
  BoothEncoderP BoothEncoderP_98 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_98_io_y),
    .io_x(BoothEncoderP_98_io_x),
    .io_p(BoothEncoderP_98_io_p)
  );
  BoothEncoderC BoothEncoderC_98 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_98_io_y),
    .io_c(BoothEncoderC_98_io_c)
  );
  BoothEncoderP BoothEncoderP_99 ( // @[CNN_CONV.scala 30:19]
    .io_y(BoothEncoderP_99_io_y),
    .io_x(BoothEncoderP_99_io_x),
    .io_p(BoothEncoderP_99_io_p)
  );
  BoothEncoderC BoothEncoderC_99 ( // @[CNN_CONV.scala 51:19]
    .io_y(BoothEncoderC_99_io_y),
    .io_c(BoothEncoderC_99_io_c)
  );
  WallaceAdder WallaceAdder ( // @[CNN_CONV.scala 213:49]
    .io_data_0(WallaceAdder_io_data_0),
    .io_data_1(WallaceAdder_io_data_1),
    .io_data_2(WallaceAdder_io_data_2),
    .io_data_3(WallaceAdder_io_data_3),
    .io_data_4(WallaceAdder_io_data_4),
    .io_data_5(WallaceAdder_io_data_5),
    .io_data_6(WallaceAdder_io_data_6),
    .io_data_7(WallaceAdder_io_data_7),
    .io_data_8(WallaceAdder_io_data_8),
    .io_data_9(WallaceAdder_io_data_9),
    .io_data_10(WallaceAdder_io_data_10),
    .io_data_11(WallaceAdder_io_data_11),
    .io_data_12(WallaceAdder_io_data_12),
    .io_data_13(WallaceAdder_io_data_13),
    .io_data_14(WallaceAdder_io_data_14),
    .io_data_15(WallaceAdder_io_data_15),
    .io_data_16(WallaceAdder_io_data_16),
    .io_data_17(WallaceAdder_io_data_17),
    .io_data_18(WallaceAdder_io_data_18),
    .io_data_19(WallaceAdder_io_data_19),
    .io_data_20(WallaceAdder_io_data_20),
    .io_data_21(WallaceAdder_io_data_21),
    .io_data_22(WallaceAdder_io_data_22),
    .io_data_23(WallaceAdder_io_data_23),
    .io_data_24(WallaceAdder_io_data_24),
    .io_cin_0(WallaceAdder_io_cin_0),
    .io_cin_1(WallaceAdder_io_cin_1),
    .io_cin_2(WallaceAdder_io_cin_2),
    .io_cin_3(WallaceAdder_io_cin_3),
    .io_cin_4(WallaceAdder_io_cin_4),
    .io_cin_5(WallaceAdder_io_cin_5),
    .io_cin_6(WallaceAdder_io_cin_6),
    .io_cin_7(WallaceAdder_io_cin_7),
    .io_cin_8(WallaceAdder_io_cin_8),
    .io_cin_9(WallaceAdder_io_cin_9),
    .io_cin_10(WallaceAdder_io_cin_10),
    .io_cin_11(WallaceAdder_io_cin_11),
    .io_cin_12(WallaceAdder_io_cin_12),
    .io_cin_13(WallaceAdder_io_cin_13),
    .io_cin_14(WallaceAdder_io_cin_14),
    .io_cin_15(WallaceAdder_io_cin_15),
    .io_cin_16(WallaceAdder_io_cin_16),
    .io_cin_17(WallaceAdder_io_cin_17),
    .io_cin_18(WallaceAdder_io_cin_18),
    .io_cin_19(WallaceAdder_io_cin_19),
    .io_cin_20(WallaceAdder_io_cin_20),
    .io_cin_21(WallaceAdder_io_cin_21),
    .io_cin_22(WallaceAdder_io_cin_22),
    .io_cin_23(WallaceAdder_io_cin_23),
    .io_cin_24(WallaceAdder_io_cin_24),
    .io_s(WallaceAdder_io_s),
    .io_c(WallaceAdder_io_c)
  );
  WallaceAdder WallaceAdder_1 ( // @[CNN_CONV.scala 213:49]
    .io_data_0(WallaceAdder_1_io_data_0),
    .io_data_1(WallaceAdder_1_io_data_1),
    .io_data_2(WallaceAdder_1_io_data_2),
    .io_data_3(WallaceAdder_1_io_data_3),
    .io_data_4(WallaceAdder_1_io_data_4),
    .io_data_5(WallaceAdder_1_io_data_5),
    .io_data_6(WallaceAdder_1_io_data_6),
    .io_data_7(WallaceAdder_1_io_data_7),
    .io_data_8(WallaceAdder_1_io_data_8),
    .io_data_9(WallaceAdder_1_io_data_9),
    .io_data_10(WallaceAdder_1_io_data_10),
    .io_data_11(WallaceAdder_1_io_data_11),
    .io_data_12(WallaceAdder_1_io_data_12),
    .io_data_13(WallaceAdder_1_io_data_13),
    .io_data_14(WallaceAdder_1_io_data_14),
    .io_data_15(WallaceAdder_1_io_data_15),
    .io_data_16(WallaceAdder_1_io_data_16),
    .io_data_17(WallaceAdder_1_io_data_17),
    .io_data_18(WallaceAdder_1_io_data_18),
    .io_data_19(WallaceAdder_1_io_data_19),
    .io_data_20(WallaceAdder_1_io_data_20),
    .io_data_21(WallaceAdder_1_io_data_21),
    .io_data_22(WallaceAdder_1_io_data_22),
    .io_data_23(WallaceAdder_1_io_data_23),
    .io_data_24(WallaceAdder_1_io_data_24),
    .io_cin_0(WallaceAdder_1_io_cin_0),
    .io_cin_1(WallaceAdder_1_io_cin_1),
    .io_cin_2(WallaceAdder_1_io_cin_2),
    .io_cin_3(WallaceAdder_1_io_cin_3),
    .io_cin_4(WallaceAdder_1_io_cin_4),
    .io_cin_5(WallaceAdder_1_io_cin_5),
    .io_cin_6(WallaceAdder_1_io_cin_6),
    .io_cin_7(WallaceAdder_1_io_cin_7),
    .io_cin_8(WallaceAdder_1_io_cin_8),
    .io_cin_9(WallaceAdder_1_io_cin_9),
    .io_cin_10(WallaceAdder_1_io_cin_10),
    .io_cin_11(WallaceAdder_1_io_cin_11),
    .io_cin_12(WallaceAdder_1_io_cin_12),
    .io_cin_13(WallaceAdder_1_io_cin_13),
    .io_cin_14(WallaceAdder_1_io_cin_14),
    .io_cin_15(WallaceAdder_1_io_cin_15),
    .io_cin_16(WallaceAdder_1_io_cin_16),
    .io_cin_17(WallaceAdder_1_io_cin_17),
    .io_cin_18(WallaceAdder_1_io_cin_18),
    .io_cin_19(WallaceAdder_1_io_cin_19),
    .io_cin_20(WallaceAdder_1_io_cin_20),
    .io_cin_21(WallaceAdder_1_io_cin_21),
    .io_cin_22(WallaceAdder_1_io_cin_22),
    .io_cin_23(WallaceAdder_1_io_cin_23),
    .io_cin_24(WallaceAdder_1_io_cin_24),
    .io_s(WallaceAdder_1_io_s),
    .io_c(WallaceAdder_1_io_c)
  );
  WallaceAdder WallaceAdder_2 ( // @[CNN_CONV.scala 213:49]
    .io_data_0(WallaceAdder_2_io_data_0),
    .io_data_1(WallaceAdder_2_io_data_1),
    .io_data_2(WallaceAdder_2_io_data_2),
    .io_data_3(WallaceAdder_2_io_data_3),
    .io_data_4(WallaceAdder_2_io_data_4),
    .io_data_5(WallaceAdder_2_io_data_5),
    .io_data_6(WallaceAdder_2_io_data_6),
    .io_data_7(WallaceAdder_2_io_data_7),
    .io_data_8(WallaceAdder_2_io_data_8),
    .io_data_9(WallaceAdder_2_io_data_9),
    .io_data_10(WallaceAdder_2_io_data_10),
    .io_data_11(WallaceAdder_2_io_data_11),
    .io_data_12(WallaceAdder_2_io_data_12),
    .io_data_13(WallaceAdder_2_io_data_13),
    .io_data_14(WallaceAdder_2_io_data_14),
    .io_data_15(WallaceAdder_2_io_data_15),
    .io_data_16(WallaceAdder_2_io_data_16),
    .io_data_17(WallaceAdder_2_io_data_17),
    .io_data_18(WallaceAdder_2_io_data_18),
    .io_data_19(WallaceAdder_2_io_data_19),
    .io_data_20(WallaceAdder_2_io_data_20),
    .io_data_21(WallaceAdder_2_io_data_21),
    .io_data_22(WallaceAdder_2_io_data_22),
    .io_data_23(WallaceAdder_2_io_data_23),
    .io_data_24(WallaceAdder_2_io_data_24),
    .io_cin_0(WallaceAdder_2_io_cin_0),
    .io_cin_1(WallaceAdder_2_io_cin_1),
    .io_cin_2(WallaceAdder_2_io_cin_2),
    .io_cin_3(WallaceAdder_2_io_cin_3),
    .io_cin_4(WallaceAdder_2_io_cin_4),
    .io_cin_5(WallaceAdder_2_io_cin_5),
    .io_cin_6(WallaceAdder_2_io_cin_6),
    .io_cin_7(WallaceAdder_2_io_cin_7),
    .io_cin_8(WallaceAdder_2_io_cin_8),
    .io_cin_9(WallaceAdder_2_io_cin_9),
    .io_cin_10(WallaceAdder_2_io_cin_10),
    .io_cin_11(WallaceAdder_2_io_cin_11),
    .io_cin_12(WallaceAdder_2_io_cin_12),
    .io_cin_13(WallaceAdder_2_io_cin_13),
    .io_cin_14(WallaceAdder_2_io_cin_14),
    .io_cin_15(WallaceAdder_2_io_cin_15),
    .io_cin_16(WallaceAdder_2_io_cin_16),
    .io_cin_17(WallaceAdder_2_io_cin_17),
    .io_cin_18(WallaceAdder_2_io_cin_18),
    .io_cin_19(WallaceAdder_2_io_cin_19),
    .io_cin_20(WallaceAdder_2_io_cin_20),
    .io_cin_21(WallaceAdder_2_io_cin_21),
    .io_cin_22(WallaceAdder_2_io_cin_22),
    .io_cin_23(WallaceAdder_2_io_cin_23),
    .io_cin_24(WallaceAdder_2_io_cin_24),
    .io_s(WallaceAdder_2_io_s),
    .io_c(WallaceAdder_2_io_c)
  );
  WallaceAdder WallaceAdder_3 ( // @[CNN_CONV.scala 213:49]
    .io_data_0(WallaceAdder_3_io_data_0),
    .io_data_1(WallaceAdder_3_io_data_1),
    .io_data_2(WallaceAdder_3_io_data_2),
    .io_data_3(WallaceAdder_3_io_data_3),
    .io_data_4(WallaceAdder_3_io_data_4),
    .io_data_5(WallaceAdder_3_io_data_5),
    .io_data_6(WallaceAdder_3_io_data_6),
    .io_data_7(WallaceAdder_3_io_data_7),
    .io_data_8(WallaceAdder_3_io_data_8),
    .io_data_9(WallaceAdder_3_io_data_9),
    .io_data_10(WallaceAdder_3_io_data_10),
    .io_data_11(WallaceAdder_3_io_data_11),
    .io_data_12(WallaceAdder_3_io_data_12),
    .io_data_13(WallaceAdder_3_io_data_13),
    .io_data_14(WallaceAdder_3_io_data_14),
    .io_data_15(WallaceAdder_3_io_data_15),
    .io_data_16(WallaceAdder_3_io_data_16),
    .io_data_17(WallaceAdder_3_io_data_17),
    .io_data_18(WallaceAdder_3_io_data_18),
    .io_data_19(WallaceAdder_3_io_data_19),
    .io_data_20(WallaceAdder_3_io_data_20),
    .io_data_21(WallaceAdder_3_io_data_21),
    .io_data_22(WallaceAdder_3_io_data_22),
    .io_data_23(WallaceAdder_3_io_data_23),
    .io_data_24(WallaceAdder_3_io_data_24),
    .io_cin_0(WallaceAdder_3_io_cin_0),
    .io_cin_1(WallaceAdder_3_io_cin_1),
    .io_cin_2(WallaceAdder_3_io_cin_2),
    .io_cin_3(WallaceAdder_3_io_cin_3),
    .io_cin_4(WallaceAdder_3_io_cin_4),
    .io_cin_5(WallaceAdder_3_io_cin_5),
    .io_cin_6(WallaceAdder_3_io_cin_6),
    .io_cin_7(WallaceAdder_3_io_cin_7),
    .io_cin_8(WallaceAdder_3_io_cin_8),
    .io_cin_9(WallaceAdder_3_io_cin_9),
    .io_cin_10(WallaceAdder_3_io_cin_10),
    .io_cin_11(WallaceAdder_3_io_cin_11),
    .io_cin_12(WallaceAdder_3_io_cin_12),
    .io_cin_13(WallaceAdder_3_io_cin_13),
    .io_cin_14(WallaceAdder_3_io_cin_14),
    .io_cin_15(WallaceAdder_3_io_cin_15),
    .io_cin_16(WallaceAdder_3_io_cin_16),
    .io_cin_17(WallaceAdder_3_io_cin_17),
    .io_cin_18(WallaceAdder_3_io_cin_18),
    .io_cin_19(WallaceAdder_3_io_cin_19),
    .io_cin_20(WallaceAdder_3_io_cin_20),
    .io_cin_21(WallaceAdder_3_io_cin_21),
    .io_cin_22(WallaceAdder_3_io_cin_22),
    .io_cin_23(WallaceAdder_3_io_cin_23),
    .io_cin_24(WallaceAdder_3_io_cin_24),
    .io_s(WallaceAdder_3_io_s),
    .io_c(WallaceAdder_3_io_c)
  );
  assign io_data_res = state ? _T_453 : res_int21; // @[CNN_CONV.scala 247:22]
  assign io_data_ok = ~stage2_valid; // @[CNN_CONV.scala 249:17]
  assign BoothEncoderP_io_y = {io_data_kernel_0[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_io_x = {16'h0,io_data_main_0}; // @[Cat.scala 30:58]
  assign BoothEncoderC_io_y = {io_data_kernel_0[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_1_io_y = {io_data_kernel_1[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_1_io_x = {16'h0,io_data_main_1}; // @[Cat.scala 30:58]
  assign BoothEncoderC_1_io_y = {io_data_kernel_1[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_2_io_y = {io_data_kernel_2[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_2_io_x = {16'h0,io_data_main_2}; // @[Cat.scala 30:58]
  assign BoothEncoderC_2_io_y = {io_data_kernel_2[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_3_io_y = {io_data_kernel_3[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_3_io_x = {16'h0,io_data_main_3}; // @[Cat.scala 30:58]
  assign BoothEncoderC_3_io_y = {io_data_kernel_3[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_4_io_y = {io_data_kernel_4[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_4_io_x = {16'h0,io_data_main_4}; // @[Cat.scala 30:58]
  assign BoothEncoderC_4_io_y = {io_data_kernel_4[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_5_io_y = {io_data_kernel_5[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_5_io_x = {16'h0,io_data_main_5}; // @[Cat.scala 30:58]
  assign BoothEncoderC_5_io_y = {io_data_kernel_5[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_6_io_y = {io_data_kernel_6[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_6_io_x = {16'h0,io_data_main_6}; // @[Cat.scala 30:58]
  assign BoothEncoderC_6_io_y = {io_data_kernel_6[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_7_io_y = {io_data_kernel_7[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_7_io_x = {16'h0,io_data_main_7}; // @[Cat.scala 30:58]
  assign BoothEncoderC_7_io_y = {io_data_kernel_7[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_8_io_y = {io_data_kernel_8[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_8_io_x = {16'h0,io_data_main_8}; // @[Cat.scala 30:58]
  assign BoothEncoderC_8_io_y = {io_data_kernel_8[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_9_io_y = {io_data_kernel_9[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_9_io_x = {16'h0,io_data_main_9}; // @[Cat.scala 30:58]
  assign BoothEncoderC_9_io_y = {io_data_kernel_9[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_10_io_y = {io_data_kernel_10[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_10_io_x = {16'h0,io_data_main_10}; // @[Cat.scala 30:58]
  assign BoothEncoderC_10_io_y = {io_data_kernel_10[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_11_io_y = {io_data_kernel_11[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_11_io_x = {16'h0,io_data_main_11}; // @[Cat.scala 30:58]
  assign BoothEncoderC_11_io_y = {io_data_kernel_11[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_12_io_y = {io_data_kernel_12[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_12_io_x = {16'h0,io_data_main_12}; // @[Cat.scala 30:58]
  assign BoothEncoderC_12_io_y = {io_data_kernel_12[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_13_io_y = {io_data_kernel_13[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_13_io_x = {16'h0,io_data_main_13}; // @[Cat.scala 30:58]
  assign BoothEncoderC_13_io_y = {io_data_kernel_13[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_14_io_y = {io_data_kernel_14[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_14_io_x = {16'h0,io_data_main_14}; // @[Cat.scala 30:58]
  assign BoothEncoderC_14_io_y = {io_data_kernel_14[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_15_io_y = {io_data_kernel_15[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_15_io_x = {16'h0,io_data_main_15}; // @[Cat.scala 30:58]
  assign BoothEncoderC_15_io_y = {io_data_kernel_15[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_16_io_y = {io_data_kernel_16[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_16_io_x = {16'h0,io_data_main_16}; // @[Cat.scala 30:58]
  assign BoothEncoderC_16_io_y = {io_data_kernel_16[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_17_io_y = {io_data_kernel_17[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_17_io_x = {16'h0,io_data_main_17}; // @[Cat.scala 30:58]
  assign BoothEncoderC_17_io_y = {io_data_kernel_17[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_18_io_y = {io_data_kernel_18[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_18_io_x = {16'h0,io_data_main_18}; // @[Cat.scala 30:58]
  assign BoothEncoderC_18_io_y = {io_data_kernel_18[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_19_io_y = {io_data_kernel_19[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_19_io_x = {16'h0,io_data_main_19}; // @[Cat.scala 30:58]
  assign BoothEncoderC_19_io_y = {io_data_kernel_19[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_20_io_y = {io_data_kernel_20[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_20_io_x = {16'h0,io_data_main_20}; // @[Cat.scala 30:58]
  assign BoothEncoderC_20_io_y = {io_data_kernel_20[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_21_io_y = {io_data_kernel_21[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_21_io_x = {16'h0,io_data_main_21}; // @[Cat.scala 30:58]
  assign BoothEncoderC_21_io_y = {io_data_kernel_21[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_22_io_y = {io_data_kernel_22[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_22_io_x = {16'h0,io_data_main_22}; // @[Cat.scala 30:58]
  assign BoothEncoderC_22_io_y = {io_data_kernel_22[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_23_io_y = {io_data_kernel_23[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_23_io_x = {16'h0,io_data_main_23}; // @[Cat.scala 30:58]
  assign BoothEncoderC_23_io_y = {io_data_kernel_23[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_24_io_y = {io_data_kernel_24[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_24_io_x = {16'h0,io_data_main_24}; // @[Cat.scala 30:58]
  assign BoothEncoderC_24_io_y = {io_data_kernel_24[1:0],1'h0}; // @[Cat.scala 30:58]
  assign BoothEncoderP_25_io_y = io_data_kernel_0[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_25_io_x = _T_127[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_25_io_y = io_data_kernel_0[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_26_io_y = io_data_kernel_1[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_26_io_x = _T_131[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_26_io_y = io_data_kernel_1[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_27_io_y = io_data_kernel_2[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_27_io_x = _T_135[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_27_io_y = io_data_kernel_2[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_28_io_y = io_data_kernel_3[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_28_io_x = _T_139[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_28_io_y = io_data_kernel_3[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_29_io_y = io_data_kernel_4[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_29_io_x = _T_143[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_29_io_y = io_data_kernel_4[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_30_io_y = io_data_kernel_5[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_30_io_x = _T_147[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_30_io_y = io_data_kernel_5[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_31_io_y = io_data_kernel_6[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_31_io_x = _T_151[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_31_io_y = io_data_kernel_6[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_32_io_y = io_data_kernel_7[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_32_io_x = _T_155[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_32_io_y = io_data_kernel_7[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_33_io_y = io_data_kernel_8[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_33_io_x = _T_159[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_33_io_y = io_data_kernel_8[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_34_io_y = io_data_kernel_9[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_34_io_x = _T_163[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_34_io_y = io_data_kernel_9[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_35_io_y = io_data_kernel_10[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_35_io_x = _T_167[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_35_io_y = io_data_kernel_10[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_36_io_y = io_data_kernel_11[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_36_io_x = _T_171[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_36_io_y = io_data_kernel_11[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_37_io_y = io_data_kernel_12[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_37_io_x = _T_175[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_37_io_y = io_data_kernel_12[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_38_io_y = io_data_kernel_13[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_38_io_x = _T_179[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_38_io_y = io_data_kernel_13[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_39_io_y = io_data_kernel_14[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_39_io_x = _T_183[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_39_io_y = io_data_kernel_14[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_40_io_y = io_data_kernel_15[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_40_io_x = _T_187[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_40_io_y = io_data_kernel_15[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_41_io_y = io_data_kernel_16[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_41_io_x = _T_191[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_41_io_y = io_data_kernel_16[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_42_io_y = io_data_kernel_17[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_42_io_x = _T_195[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_42_io_y = io_data_kernel_17[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_43_io_y = io_data_kernel_18[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_43_io_x = _T_199[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_43_io_y = io_data_kernel_18[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_44_io_y = io_data_kernel_19[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_44_io_x = _T_203[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_44_io_y = io_data_kernel_19[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_45_io_y = io_data_kernel_20[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_45_io_x = _T_207[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_45_io_y = io_data_kernel_20[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_46_io_y = io_data_kernel_21[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_46_io_x = _T_211[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_46_io_y = io_data_kernel_21[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_47_io_y = io_data_kernel_22[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_47_io_x = _T_215[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_47_io_y = io_data_kernel_22[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_48_io_y = io_data_kernel_23[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_48_io_x = _T_219[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_48_io_y = io_data_kernel_23[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_49_io_y = io_data_kernel_24[3:1]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_49_io_x = _T_223[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_49_io_y = io_data_kernel_24[3:1]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_50_io_y = io_data_kernel_0[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_50_io_x = _T_227[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_50_io_y = io_data_kernel_0[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_51_io_y = io_data_kernel_1[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_51_io_x = _T_231[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_51_io_y = io_data_kernel_1[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_52_io_y = io_data_kernel_2[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_52_io_x = _T_235[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_52_io_y = io_data_kernel_2[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_53_io_y = io_data_kernel_3[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_53_io_x = _T_239[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_53_io_y = io_data_kernel_3[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_54_io_y = io_data_kernel_4[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_54_io_x = _T_243[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_54_io_y = io_data_kernel_4[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_55_io_y = io_data_kernel_5[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_55_io_x = _T_247[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_55_io_y = io_data_kernel_5[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_56_io_y = io_data_kernel_6[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_56_io_x = _T_251[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_56_io_y = io_data_kernel_6[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_57_io_y = io_data_kernel_7[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_57_io_x = _T_255[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_57_io_y = io_data_kernel_7[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_58_io_y = io_data_kernel_8[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_58_io_x = _T_259[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_58_io_y = io_data_kernel_8[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_59_io_y = io_data_kernel_9[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_59_io_x = _T_263[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_59_io_y = io_data_kernel_9[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_60_io_y = io_data_kernel_10[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_60_io_x = _T_267[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_60_io_y = io_data_kernel_10[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_61_io_y = io_data_kernel_11[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_61_io_x = _T_271[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_61_io_y = io_data_kernel_11[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_62_io_y = io_data_kernel_12[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_62_io_x = _T_275[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_62_io_y = io_data_kernel_12[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_63_io_y = io_data_kernel_13[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_63_io_x = _T_279[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_63_io_y = io_data_kernel_13[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_64_io_y = io_data_kernel_14[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_64_io_x = _T_283[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_64_io_y = io_data_kernel_14[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_65_io_y = io_data_kernel_15[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_65_io_x = _T_287[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_65_io_y = io_data_kernel_15[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_66_io_y = io_data_kernel_16[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_66_io_x = _T_291[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_66_io_y = io_data_kernel_16[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_67_io_y = io_data_kernel_17[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_67_io_x = _T_295[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_67_io_y = io_data_kernel_17[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_68_io_y = io_data_kernel_18[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_68_io_x = _T_299[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_68_io_y = io_data_kernel_18[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_69_io_y = io_data_kernel_19[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_69_io_x = _T_303[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_69_io_y = io_data_kernel_19[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_70_io_y = io_data_kernel_20[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_70_io_x = _T_307[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_70_io_y = io_data_kernel_20[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_71_io_y = io_data_kernel_21[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_71_io_x = _T_311[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_71_io_y = io_data_kernel_21[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_72_io_y = io_data_kernel_22[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_72_io_x = _T_315[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_72_io_y = io_data_kernel_22[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_73_io_y = io_data_kernel_23[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_73_io_x = _T_319[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_73_io_y = io_data_kernel_23[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_74_io_y = io_data_kernel_24[5:3]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_74_io_x = _T_323[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_74_io_y = io_data_kernel_24[5:3]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_75_io_y = io_data_kernel_0[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_75_io_x = _T_327[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_75_io_y = io_data_kernel_0[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_76_io_y = io_data_kernel_1[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_76_io_x = _T_331[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_76_io_y = io_data_kernel_1[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_77_io_y = io_data_kernel_2[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_77_io_x = _T_335[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_77_io_y = io_data_kernel_2[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_78_io_y = io_data_kernel_3[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_78_io_x = _T_339[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_78_io_y = io_data_kernel_3[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_79_io_y = io_data_kernel_4[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_79_io_x = _T_343[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_79_io_y = io_data_kernel_4[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_80_io_y = io_data_kernel_5[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_80_io_x = _T_347[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_80_io_y = io_data_kernel_5[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_81_io_y = io_data_kernel_6[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_81_io_x = _T_351[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_81_io_y = io_data_kernel_6[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_82_io_y = io_data_kernel_7[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_82_io_x = _T_355[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_82_io_y = io_data_kernel_7[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_83_io_y = io_data_kernel_8[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_83_io_x = _T_359[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_83_io_y = io_data_kernel_8[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_84_io_y = io_data_kernel_9[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_84_io_x = _T_363[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_84_io_y = io_data_kernel_9[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_85_io_y = io_data_kernel_10[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_85_io_x = _T_367[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_85_io_y = io_data_kernel_10[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_86_io_y = io_data_kernel_11[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_86_io_x = _T_371[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_86_io_y = io_data_kernel_11[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_87_io_y = io_data_kernel_12[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_87_io_x = _T_375[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_87_io_y = io_data_kernel_12[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_88_io_y = io_data_kernel_13[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_88_io_x = _T_379[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_88_io_y = io_data_kernel_13[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_89_io_y = io_data_kernel_14[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_89_io_x = _T_383[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_89_io_y = io_data_kernel_14[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_90_io_y = io_data_kernel_15[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_90_io_x = _T_387[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_90_io_y = io_data_kernel_15[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_91_io_y = io_data_kernel_16[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_91_io_x = _T_391[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_91_io_y = io_data_kernel_16[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_92_io_y = io_data_kernel_17[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_92_io_x = _T_395[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_92_io_y = io_data_kernel_17[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_93_io_y = io_data_kernel_18[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_93_io_x = _T_399[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_93_io_y = io_data_kernel_18[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_94_io_y = io_data_kernel_19[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_94_io_x = _T_403[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_94_io_y = io_data_kernel_19[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_95_io_y = io_data_kernel_20[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_95_io_x = _T_407[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_95_io_y = io_data_kernel_20[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_96_io_y = io_data_kernel_21[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_96_io_x = _T_411[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_96_io_y = io_data_kernel_21[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_97_io_y = io_data_kernel_22[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_97_io_x = _T_415[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_97_io_y = io_data_kernel_22[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_98_io_y = io_data_kernel_23[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_98_io_x = _T_419[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_98_io_y = io_data_kernel_23[7:5]; // @[CNN_CONV.scala 207:58]
  assign BoothEncoderP_99_io_y = io_data_kernel_24[7:5]; // @[CNN_CONV.scala 206:58]
  assign BoothEncoderP_99_io_x = _T_423[31:0]; // @[CNN_CONV.scala 32:12]
  assign BoothEncoderC_99_io_y = io_data_kernel_24[7:5]; // @[CNN_CONV.scala 207:58]
  assign WallaceAdder_io_data_0 = BoothEncoderP_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_1 = BoothEncoderP_1_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_2 = BoothEncoderP_2_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_3 = BoothEncoderP_3_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_4 = BoothEncoderP_4_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_5 = BoothEncoderP_5_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_6 = BoothEncoderP_6_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_7 = BoothEncoderP_7_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_8 = BoothEncoderP_8_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_9 = BoothEncoderP_9_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_10 = BoothEncoderP_10_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_11 = BoothEncoderP_11_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_12 = BoothEncoderP_12_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_13 = BoothEncoderP_13_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_14 = BoothEncoderP_14_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_15 = BoothEncoderP_15_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_16 = BoothEncoderP_16_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_17 = BoothEncoderP_17_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_18 = BoothEncoderP_18_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_19 = BoothEncoderP_19_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_20 = BoothEncoderP_20_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_21 = BoothEncoderP_21_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_22 = BoothEncoderP_22_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_23 = BoothEncoderP_23_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_data_24 = BoothEncoderP_24_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_io_cin_0 = BoothEncoderC_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_1 = BoothEncoderC_1_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_2 = BoothEncoderC_2_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_3 = BoothEncoderC_3_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_4 = BoothEncoderC_4_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_5 = BoothEncoderC_5_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_6 = BoothEncoderC_6_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_7 = BoothEncoderC_7_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_8 = BoothEncoderC_8_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_9 = BoothEncoderC_9_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_10 = BoothEncoderC_10_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_11 = BoothEncoderC_11_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_12 = BoothEncoderC_12_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_13 = BoothEncoderC_13_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_14 = BoothEncoderC_14_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_15 = BoothEncoderC_15_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_16 = BoothEncoderC_16_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_17 = BoothEncoderC_17_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_18 = BoothEncoderC_18_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_19 = BoothEncoderC_19_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_20 = BoothEncoderC_20_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_21 = BoothEncoderC_21_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_22 = BoothEncoderC_22_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_23 = BoothEncoderC_23_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_io_cin_24 = BoothEncoderC_24_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_data_0 = BoothEncoderP_25_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_1 = BoothEncoderP_26_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_2 = BoothEncoderP_27_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_3 = BoothEncoderP_28_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_4 = BoothEncoderP_29_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_5 = BoothEncoderP_30_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_6 = BoothEncoderP_31_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_7 = BoothEncoderP_32_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_8 = BoothEncoderP_33_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_9 = BoothEncoderP_34_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_10 = BoothEncoderP_35_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_11 = BoothEncoderP_36_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_12 = BoothEncoderP_37_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_13 = BoothEncoderP_38_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_14 = BoothEncoderP_39_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_15 = BoothEncoderP_40_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_16 = BoothEncoderP_41_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_17 = BoothEncoderP_42_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_18 = BoothEncoderP_43_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_19 = BoothEncoderP_44_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_20 = BoothEncoderP_45_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_21 = BoothEncoderP_46_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_22 = BoothEncoderP_47_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_23 = BoothEncoderP_48_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_data_24 = BoothEncoderP_49_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_1_io_cin_0 = BoothEncoderC_25_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_1 = BoothEncoderC_26_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_2 = BoothEncoderC_27_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_3 = BoothEncoderC_28_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_4 = BoothEncoderC_29_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_5 = BoothEncoderC_30_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_6 = BoothEncoderC_31_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_7 = BoothEncoderC_32_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_8 = BoothEncoderC_33_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_9 = BoothEncoderC_34_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_10 = BoothEncoderC_35_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_11 = BoothEncoderC_36_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_12 = BoothEncoderC_37_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_13 = BoothEncoderC_38_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_14 = BoothEncoderC_39_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_15 = BoothEncoderC_40_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_16 = BoothEncoderC_41_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_17 = BoothEncoderC_42_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_18 = BoothEncoderC_43_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_19 = BoothEncoderC_44_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_20 = BoothEncoderC_45_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_21 = BoothEncoderC_46_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_22 = BoothEncoderC_47_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_23 = BoothEncoderC_48_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_1_io_cin_24 = BoothEncoderC_49_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_data_0 = BoothEncoderP_50_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_1 = BoothEncoderP_51_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_2 = BoothEncoderP_52_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_3 = BoothEncoderP_53_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_4 = BoothEncoderP_54_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_5 = BoothEncoderP_55_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_6 = BoothEncoderP_56_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_7 = BoothEncoderP_57_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_8 = BoothEncoderP_58_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_9 = BoothEncoderP_59_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_10 = BoothEncoderP_60_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_11 = BoothEncoderP_61_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_12 = BoothEncoderP_62_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_13 = BoothEncoderP_63_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_14 = BoothEncoderP_64_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_15 = BoothEncoderP_65_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_16 = BoothEncoderP_66_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_17 = BoothEncoderP_67_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_18 = BoothEncoderP_68_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_19 = BoothEncoderP_69_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_20 = BoothEncoderP_70_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_21 = BoothEncoderP_71_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_22 = BoothEncoderP_72_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_23 = BoothEncoderP_73_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_data_24 = BoothEncoderP_74_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_2_io_cin_0 = BoothEncoderC_50_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_1 = BoothEncoderC_51_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_2 = BoothEncoderC_52_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_3 = BoothEncoderC_53_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_4 = BoothEncoderC_54_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_5 = BoothEncoderC_55_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_6 = BoothEncoderC_56_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_7 = BoothEncoderC_57_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_8 = BoothEncoderC_58_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_9 = BoothEncoderC_59_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_10 = BoothEncoderC_60_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_11 = BoothEncoderC_61_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_12 = BoothEncoderC_62_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_13 = BoothEncoderC_63_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_14 = BoothEncoderC_64_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_15 = BoothEncoderC_65_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_16 = BoothEncoderC_66_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_17 = BoothEncoderC_67_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_18 = BoothEncoderC_68_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_19 = BoothEncoderC_69_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_20 = BoothEncoderC_70_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_21 = BoothEncoderC_71_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_22 = BoothEncoderC_72_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_23 = BoothEncoderC_73_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_2_io_cin_24 = BoothEncoderC_74_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_data_0 = BoothEncoderP_75_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_1 = BoothEncoderP_76_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_2 = BoothEncoderP_77_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_3 = BoothEncoderP_78_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_4 = BoothEncoderP_79_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_5 = BoothEncoderP_80_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_6 = BoothEncoderP_81_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_7 = BoothEncoderP_82_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_8 = BoothEncoderP_83_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_9 = BoothEncoderP_84_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_10 = BoothEncoderP_85_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_11 = BoothEncoderP_86_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_12 = BoothEncoderP_87_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_13 = BoothEncoderP_88_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_14 = BoothEncoderP_89_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_15 = BoothEncoderP_90_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_16 = BoothEncoderP_91_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_17 = BoothEncoderP_92_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_18 = BoothEncoderP_93_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_19 = BoothEncoderP_94_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_20 = BoothEncoderP_95_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_21 = BoothEncoderP_96_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_22 = BoothEncoderP_97_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_23 = BoothEncoderP_98_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_data_24 = BoothEncoderP_99_io_p; // @[CNN_CONV.scala 213:30 217:27]
  assign WallaceAdder_3_io_cin_0 = BoothEncoderC_75_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_1 = BoothEncoderC_76_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_2 = BoothEncoderC_77_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_3 = BoothEncoderC_78_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_4 = BoothEncoderC_79_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_5 = BoothEncoderC_80_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_6 = BoothEncoderC_81_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_7 = BoothEncoderC_82_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_8 = BoothEncoderC_83_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_9 = BoothEncoderC_84_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_10 = BoothEncoderC_85_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_11 = BoothEncoderC_86_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_12 = BoothEncoderC_87_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_13 = BoothEncoderC_88_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_14 = BoothEncoderC_89_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_15 = BoothEncoderC_90_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_16 = BoothEncoderC_91_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_17 = BoothEncoderC_92_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_18 = BoothEncoderC_93_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_19 = BoothEncoderC_94_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_20 = BoothEncoderC_95_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_21 = BoothEncoderC_96_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_22 = BoothEncoderC_97_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_23 = BoothEncoderC_98_io_c; // @[CNN_CONV.scala 213:30 218:27]
  assign WallaceAdder_3_io_cin_24 = BoothEncoderC_99_io_c; // @[CNN_CONV.scala 213:30 218:27]
  always @(posedge clock) begin
    if (reset) begin // @[CNN_CONV.scala 228:22]
      state <= 1'h0; // @[CNN_CONV.scala 228:22]
    end else if (_T_426) begin // @[CNN_CONV.scala 230:18]
      state <= _GEN_0;
    end else if (state) begin // @[CNN_CONV.scala 230:18]
      state <= 1'h0; // @[CNN_CONV.scala 235:13]
    end
    if (reset) begin // @[CNN_CONV.scala 238:26]
      out_s_reg_0 <= 32'h0; // @[CNN_CONV.scala 238:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 240:23]
      out_s_reg_0 <= wallace_adder_0_s; // @[CNN_CONV.scala 240:35]
    end
    if (reset) begin // @[CNN_CONV.scala 238:26]
      out_s_reg_1 <= 32'h0; // @[CNN_CONV.scala 238:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 240:23]
      out_s_reg_1 <= wallace_adder_1_s; // @[CNN_CONV.scala 240:35]
    end
    if (reset) begin // @[CNN_CONV.scala 238:26]
      out_s_reg_2 <= 32'h0; // @[CNN_CONV.scala 238:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 240:23]
      out_s_reg_2 <= wallace_adder_2_s; // @[CNN_CONV.scala 240:35]
    end
    if (reset) begin // @[CNN_CONV.scala 238:26]
      out_s_reg_3 <= 32'h0; // @[CNN_CONV.scala 238:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 240:23]
      out_s_reg_3 <= wallace_adder_3_s; // @[CNN_CONV.scala 240:35]
    end
    if (reset) begin // @[CNN_CONV.scala 239:26]
      out_c_reg_0 <= 32'h0; // @[CNN_CONV.scala 239:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 241:23]
      out_c_reg_0 <= wallace_adder_0_c; // @[CNN_CONV.scala 241:35]
    end
    if (reset) begin // @[CNN_CONV.scala 239:26]
      out_c_reg_1 <= 32'h0; // @[CNN_CONV.scala 239:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 241:23]
      out_c_reg_1 <= wallace_adder_1_c; // @[CNN_CONV.scala 241:35]
    end
    if (reset) begin // @[CNN_CONV.scala 239:26]
      out_c_reg_2 <= 32'h0; // @[CNN_CONV.scala 239:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 241:23]
      out_c_reg_2 <= wallace_adder_2_c; // @[CNN_CONV.scala 241:35]
    end
    if (reset) begin // @[CNN_CONV.scala 239:26]
      out_c_reg_3 <= 32'h0; // @[CNN_CONV.scala 239:26]
    end else if (stage2_valid) begin // @[CNN_CONV.scala 241:23]
      out_c_reg_3 <= wallace_adder_3_c; // @[CNN_CONV.scala 241:35]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_s_reg_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  out_s_reg_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  out_s_reg_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  out_s_reg_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  out_c_reg_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  out_c_reg_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  out_c_reg_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  out_c_reg_3 = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CNNConv(
  input         clock,
  input         reset,
  input         io_conv_valid,
  input  [15:0] io_data_main_0,
  input  [15:0] io_data_main_1,
  input  [15:0] io_data_main_2,
  input  [15:0] io_data_main_3,
  input  [15:0] io_data_main_4,
  input  [15:0] io_data_main_5,
  input  [15:0] io_data_main_6,
  input  [15:0] io_data_main_7,
  input  [15:0] io_data_main_8,
  input  [15:0] io_data_main_9,
  input  [15:0] io_data_main_10,
  input  [15:0] io_data_main_11,
  input  [15:0] io_data_main_12,
  input  [15:0] io_data_main_13,
  input  [15:0] io_data_main_14,
  input  [15:0] io_data_main_15,
  input  [15:0] io_data_main_16,
  input  [15:0] io_data_main_17,
  input  [15:0] io_data_main_18,
  input  [15:0] io_data_main_19,
  input  [15:0] io_data_main_20,
  input  [15:0] io_data_main_21,
  input  [15:0] io_data_main_22,
  input  [15:0] io_data_main_23,
  input  [15:0] io_data_main_24,
  input  [7:0]  io_data_kernel_0,
  input  [7:0]  io_data_kernel_1,
  input  [7:0]  io_data_kernel_2,
  input  [7:0]  io_data_kernel_3,
  input  [7:0]  io_data_kernel_4,
  input  [7:0]  io_data_kernel_5,
  input  [7:0]  io_data_kernel_6,
  input  [7:0]  io_data_kernel_7,
  input  [7:0]  io_data_kernel_8,
  input  [7:0]  io_data_kernel_9,
  input  [7:0]  io_data_kernel_10,
  input  [7:0]  io_data_kernel_11,
  input  [7:0]  io_data_kernel_12,
  input  [7:0]  io_data_kernel_13,
  input  [7:0]  io_data_kernel_14,
  input  [7:0]  io_data_kernel_15,
  input  [7:0]  io_data_kernel_16,
  input  [7:0]  io_data_kernel_17,
  input  [7:0]  io_data_kernel_18,
  input  [7:0]  io_data_kernel_19,
  input  [7:0]  io_data_kernel_20,
  input  [7:0]  io_data_kernel_21,
  input  [7:0]  io_data_kernel_22,
  input  [7:0]  io_data_kernel_23,
  input  [7:0]  io_data_kernel_24,
  input  [3:0]  io_data_kernel_vwidth,
  output [63:0] io_conv_res,
  output        io_conv_ok
);
  wire  conv_mdu_clock; // @[CNN_CONV.scala 271:24]
  wire  conv_mdu_reset; // @[CNN_CONV.scala 271:24]
  wire  conv_mdu_io_conv_valid; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_0; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_1; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_2; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_3; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_4; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_5; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_6; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_7; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_8; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_9; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_10; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_11; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_12; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_13; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_14; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_15; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_16; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_17; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_18; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_19; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_20; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_21; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_22; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_23; // @[CNN_CONV.scala 271:24]
  wire [15:0] conv_mdu_io_data_main_24; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_0; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_1; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_2; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_3; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_4; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_5; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_6; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_7; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_8; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_9; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_10; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_11; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_12; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_13; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_14; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_15; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_16; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_17; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_18; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_19; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_20; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_21; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_22; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_23; // @[CNN_CONV.scala 271:24]
  wire [7:0] conv_mdu_io_data_kernel_24; // @[CNN_CONV.scala 271:24]
  wire [3:0] conv_mdu_io_data_kernel_vwidth; // @[CNN_CONV.scala 271:24]
  wire [31:0] conv_mdu_io_data_res; // @[CNN_CONV.scala 271:24]
  wire  conv_mdu_io_data_ok; // @[CNN_CONV.scala 271:24]
  CNNConvSub25 conv_mdu ( // @[CNN_CONV.scala 271:24]
    .clock(conv_mdu_clock),
    .reset(conv_mdu_reset),
    .io_conv_valid(conv_mdu_io_conv_valid),
    .io_data_main_0(conv_mdu_io_data_main_0),
    .io_data_main_1(conv_mdu_io_data_main_1),
    .io_data_main_2(conv_mdu_io_data_main_2),
    .io_data_main_3(conv_mdu_io_data_main_3),
    .io_data_main_4(conv_mdu_io_data_main_4),
    .io_data_main_5(conv_mdu_io_data_main_5),
    .io_data_main_6(conv_mdu_io_data_main_6),
    .io_data_main_7(conv_mdu_io_data_main_7),
    .io_data_main_8(conv_mdu_io_data_main_8),
    .io_data_main_9(conv_mdu_io_data_main_9),
    .io_data_main_10(conv_mdu_io_data_main_10),
    .io_data_main_11(conv_mdu_io_data_main_11),
    .io_data_main_12(conv_mdu_io_data_main_12),
    .io_data_main_13(conv_mdu_io_data_main_13),
    .io_data_main_14(conv_mdu_io_data_main_14),
    .io_data_main_15(conv_mdu_io_data_main_15),
    .io_data_main_16(conv_mdu_io_data_main_16),
    .io_data_main_17(conv_mdu_io_data_main_17),
    .io_data_main_18(conv_mdu_io_data_main_18),
    .io_data_main_19(conv_mdu_io_data_main_19),
    .io_data_main_20(conv_mdu_io_data_main_20),
    .io_data_main_21(conv_mdu_io_data_main_21),
    .io_data_main_22(conv_mdu_io_data_main_22),
    .io_data_main_23(conv_mdu_io_data_main_23),
    .io_data_main_24(conv_mdu_io_data_main_24),
    .io_data_kernel_0(conv_mdu_io_data_kernel_0),
    .io_data_kernel_1(conv_mdu_io_data_kernel_1),
    .io_data_kernel_2(conv_mdu_io_data_kernel_2),
    .io_data_kernel_3(conv_mdu_io_data_kernel_3),
    .io_data_kernel_4(conv_mdu_io_data_kernel_4),
    .io_data_kernel_5(conv_mdu_io_data_kernel_5),
    .io_data_kernel_6(conv_mdu_io_data_kernel_6),
    .io_data_kernel_7(conv_mdu_io_data_kernel_7),
    .io_data_kernel_8(conv_mdu_io_data_kernel_8),
    .io_data_kernel_9(conv_mdu_io_data_kernel_9),
    .io_data_kernel_10(conv_mdu_io_data_kernel_10),
    .io_data_kernel_11(conv_mdu_io_data_kernel_11),
    .io_data_kernel_12(conv_mdu_io_data_kernel_12),
    .io_data_kernel_13(conv_mdu_io_data_kernel_13),
    .io_data_kernel_14(conv_mdu_io_data_kernel_14),
    .io_data_kernel_15(conv_mdu_io_data_kernel_15),
    .io_data_kernel_16(conv_mdu_io_data_kernel_16),
    .io_data_kernel_17(conv_mdu_io_data_kernel_17),
    .io_data_kernel_18(conv_mdu_io_data_kernel_18),
    .io_data_kernel_19(conv_mdu_io_data_kernel_19),
    .io_data_kernel_20(conv_mdu_io_data_kernel_20),
    .io_data_kernel_21(conv_mdu_io_data_kernel_21),
    .io_data_kernel_22(conv_mdu_io_data_kernel_22),
    .io_data_kernel_23(conv_mdu_io_data_kernel_23),
    .io_data_kernel_24(conv_mdu_io_data_kernel_24),
    .io_data_kernel_vwidth(conv_mdu_io_data_kernel_vwidth),
    .io_data_res(conv_mdu_io_data_res),
    .io_data_ok(conv_mdu_io_data_ok)
  );
  assign io_conv_res = {32'h0,conv_mdu_io_data_res}; // @[Cat.scala 30:58]
  assign io_conv_ok = conv_mdu_io_data_ok; // @[CNN_CONV.scala 288:14]
  assign conv_mdu_clock = clock;
  assign conv_mdu_reset = reset;
  assign conv_mdu_io_conv_valid = io_conv_valid; // @[CNN_CONV.scala 272:26]
  assign conv_mdu_io_data_main_0 = io_data_main_0; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_1 = io_data_main_1; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_2 = io_data_main_2; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_3 = io_data_main_3; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_4 = io_data_main_4; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_5 = io_data_main_5; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_6 = io_data_main_6; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_7 = io_data_main_7; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_8 = io_data_main_8; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_9 = io_data_main_9; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_10 = io_data_main_10; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_11 = io_data_main_11; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_12 = io_data_main_12; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_13 = io_data_main_13; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_14 = io_data_main_14; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_15 = io_data_main_15; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_16 = io_data_main_16; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_17 = io_data_main_17; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_18 = io_data_main_18; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_19 = io_data_main_19; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_20 = io_data_main_20; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_21 = io_data_main_21; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_22 = io_data_main_22; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_23 = io_data_main_23; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_main_24 = io_data_main_24; // @[CNN_CONV.scala 273:25]
  assign conv_mdu_io_data_kernel_0 = io_data_kernel_0; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_1 = io_data_kernel_1; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_2 = io_data_kernel_2; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_3 = io_data_kernel_3; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_4 = io_data_kernel_4; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_5 = io_data_kernel_5; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_6 = io_data_kernel_6; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_7 = io_data_kernel_7; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_8 = io_data_kernel_8; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_9 = io_data_kernel_9; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_10 = io_data_kernel_10; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_11 = io_data_kernel_11; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_12 = io_data_kernel_12; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_13 = io_data_kernel_13; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_14 = io_data_kernel_14; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_15 = io_data_kernel_15; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_16 = io_data_kernel_16; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_17 = io_data_kernel_17; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_18 = io_data_kernel_18; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_19 = io_data_kernel_19; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_20 = io_data_kernel_20; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_21 = io_data_kernel_21; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_22 = io_data_kernel_22; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_23 = io_data_kernel_23; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_24 = io_data_kernel_24; // @[CNN_CONV.scala 274:27]
  assign conv_mdu_io_data_kernel_vwidth = io_data_kernel_vwidth; // @[CNN_CONV.scala 275:34]
endmodule
module CNNPoolMax(
  input  [15:0] io_data_main_0,
  input  [15:0] io_data_main_1,
  input  [15:0] io_data_main_2,
  input  [15:0] io_data_main_3,
  input  [15:0] io_data_main_4,
  input  [15:0] io_data_main_5,
  input  [15:0] io_data_main_6,
  input  [15:0] io_data_main_7,
  input  [15:0] io_data_main_8,
  input  [15:0] io_data_main_9,
  input  [15:0] io_data_main_10,
  input  [15:0] io_data_main_11,
  input  [15:0] io_data_main_12,
  input  [15:0] io_data_main_13,
  input  [15:0] io_data_main_14,
  input  [15:0] io_data_main_15,
  input  [15:0] io_data_main_16,
  input  [15:0] io_data_main_17,
  input  [15:0] io_data_main_18,
  input  [15:0] io_data_main_19,
  input  [15:0] io_data_main_20,
  input  [15:0] io_data_main_21,
  input  [15:0] io_data_main_22,
  input  [15:0] io_data_main_23,
  input  [15:0] io_data_main_24,
  output [15:0] io_data_res
);
  wire [15:0] _T_1 = io_data_main_0 >= io_data_main_1 ? io_data_main_0 : io_data_main_1; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_3 = _T_1 >= io_data_main_2 ? _T_1 : io_data_main_2; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_5 = _T_3 >= io_data_main_3 ? _T_3 : io_data_main_3; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_7 = _T_5 >= io_data_main_4 ? _T_5 : io_data_main_4; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_9 = _T_7 >= io_data_main_5 ? _T_7 : io_data_main_5; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_11 = _T_9 >= io_data_main_6 ? _T_9 : io_data_main_6; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_13 = _T_11 >= io_data_main_7 ? _T_11 : io_data_main_7; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_15 = _T_13 >= io_data_main_8 ? _T_13 : io_data_main_8; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_17 = _T_15 >= io_data_main_9 ? _T_15 : io_data_main_9; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_19 = _T_17 >= io_data_main_10 ? _T_17 : io_data_main_10; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_21 = _T_19 >= io_data_main_11 ? _T_19 : io_data_main_11; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_23 = _T_21 >= io_data_main_12 ? _T_21 : io_data_main_12; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_25 = _T_23 >= io_data_main_13 ? _T_23 : io_data_main_13; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_27 = _T_25 >= io_data_main_14 ? _T_25 : io_data_main_14; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_29 = _T_27 >= io_data_main_15 ? _T_27 : io_data_main_15; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_31 = _T_29 >= io_data_main_16 ? _T_29 : io_data_main_16; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_33 = _T_31 >= io_data_main_17 ? _T_31 : io_data_main_17; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_35 = _T_33 >= io_data_main_18 ? _T_33 : io_data_main_18; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_37 = _T_35 >= io_data_main_19 ? _T_35 : io_data_main_19; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_39 = _T_37 >= io_data_main_20 ? _T_37 : io_data_main_20; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_41 = _T_39 >= io_data_main_21 ? _T_39 : io_data_main_21; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_43 = _T_41 >= io_data_main_22 ? _T_41 : io_data_main_22; // @[CNN_POOL.scala 15:52]
  wire [15:0] _T_45 = _T_43 >= io_data_main_23 ? _T_43 : io_data_main_23; // @[CNN_POOL.scala 15:52]
  assign io_data_res = _T_45 >= io_data_main_24 ? _T_45 : io_data_main_24; // @[CNN_POOL.scala 15:52]
endmodule
module CNNPoolAvg(
  input  [3:0]  io_k,
  input  [15:0] io_data_main_0,
  input  [15:0] io_data_main_1,
  input  [15:0] io_data_main_2,
  input  [15:0] io_data_main_3,
  input  [15:0] io_data_main_4,
  input  [15:0] io_data_main_5,
  input  [15:0] io_data_main_6,
  input  [15:0] io_data_main_7,
  input  [15:0] io_data_main_8,
  input  [15:0] io_data_main_9,
  input  [15:0] io_data_main_10,
  input  [15:0] io_data_main_11,
  input  [15:0] io_data_main_12,
  input  [15:0] io_data_main_13,
  input  [15:0] io_data_main_14,
  input  [15:0] io_data_main_15,
  input  [15:0] io_data_main_16,
  input  [15:0] io_data_main_17,
  input  [15:0] io_data_main_18,
  input  [15:0] io_data_main_19,
  input  [15:0] io_data_main_20,
  input  [15:0] io_data_main_21,
  input  [15:0] io_data_main_22,
  input  [15:0] io_data_main_23,
  input  [15:0] io_data_main_24,
  output [15:0] io_data_res
);
  wire [16:0] _T = io_data_main_0 + io_data_main_1; // @[CNN_POOL.scala 26:32]
  wire [16:0] _GEN_0 = {{1'd0}, io_data_main_2}; // @[CNN_POOL.scala 26:32]
  wire [17:0] _T_1 = _T + _GEN_0; // @[CNN_POOL.scala 26:32]
  wire [17:0] _GEN_1 = {{2'd0}, io_data_main_3}; // @[CNN_POOL.scala 26:32]
  wire [18:0] _T_2 = _T_1 + _GEN_1; // @[CNN_POOL.scala 26:32]
  wire [18:0] _GEN_2 = {{3'd0}, io_data_main_4}; // @[CNN_POOL.scala 26:32]
  wire [19:0] _T_3 = _T_2 + _GEN_2; // @[CNN_POOL.scala 26:32]
  wire [19:0] _GEN_3 = {{4'd0}, io_data_main_5}; // @[CNN_POOL.scala 26:32]
  wire [20:0] _T_4 = _T_3 + _GEN_3; // @[CNN_POOL.scala 26:32]
  wire [20:0] _GEN_4 = {{5'd0}, io_data_main_6}; // @[CNN_POOL.scala 26:32]
  wire [21:0] _T_5 = _T_4 + _GEN_4; // @[CNN_POOL.scala 26:32]
  wire [21:0] _GEN_5 = {{6'd0}, io_data_main_7}; // @[CNN_POOL.scala 26:32]
  wire [22:0] _T_6 = _T_5 + _GEN_5; // @[CNN_POOL.scala 26:32]
  wire [22:0] _GEN_6 = {{7'd0}, io_data_main_8}; // @[CNN_POOL.scala 26:32]
  wire [23:0] _T_7 = _T_6 + _GEN_6; // @[CNN_POOL.scala 26:32]
  wire [23:0] _GEN_7 = {{8'd0}, io_data_main_9}; // @[CNN_POOL.scala 26:32]
  wire [24:0] _T_8 = _T_7 + _GEN_7; // @[CNN_POOL.scala 26:32]
  wire [24:0] _GEN_8 = {{9'd0}, io_data_main_10}; // @[CNN_POOL.scala 26:32]
  wire [25:0] _T_9 = _T_8 + _GEN_8; // @[CNN_POOL.scala 26:32]
  wire [25:0] _GEN_9 = {{10'd0}, io_data_main_11}; // @[CNN_POOL.scala 26:32]
  wire [26:0] _T_10 = _T_9 + _GEN_9; // @[CNN_POOL.scala 26:32]
  wire [26:0] _GEN_10 = {{11'd0}, io_data_main_12}; // @[CNN_POOL.scala 26:32]
  wire [27:0] _T_11 = _T_10 + _GEN_10; // @[CNN_POOL.scala 26:32]
  wire [27:0] _GEN_11 = {{12'd0}, io_data_main_13}; // @[CNN_POOL.scala 26:32]
  wire [28:0] _T_12 = _T_11 + _GEN_11; // @[CNN_POOL.scala 26:32]
  wire [28:0] _GEN_12 = {{13'd0}, io_data_main_14}; // @[CNN_POOL.scala 26:32]
  wire [29:0] _T_13 = _T_12 + _GEN_12; // @[CNN_POOL.scala 26:32]
  wire [29:0] _GEN_13 = {{14'd0}, io_data_main_15}; // @[CNN_POOL.scala 26:32]
  wire [30:0] _T_14 = _T_13 + _GEN_13; // @[CNN_POOL.scala 26:32]
  wire [30:0] _GEN_14 = {{15'd0}, io_data_main_16}; // @[CNN_POOL.scala 26:32]
  wire [31:0] _T_15 = _T_14 + _GEN_14; // @[CNN_POOL.scala 26:32]
  wire [31:0] _GEN_15 = {{16'd0}, io_data_main_17}; // @[CNN_POOL.scala 26:32]
  wire [32:0] _T_16 = _T_15 + _GEN_15; // @[CNN_POOL.scala 26:32]
  wire [32:0] _GEN_16 = {{17'd0}, io_data_main_18}; // @[CNN_POOL.scala 26:32]
  wire [33:0] _T_17 = _T_16 + _GEN_16; // @[CNN_POOL.scala 26:32]
  wire [33:0] _GEN_17 = {{18'd0}, io_data_main_19}; // @[CNN_POOL.scala 26:32]
  wire [34:0] _T_18 = _T_17 + _GEN_17; // @[CNN_POOL.scala 26:32]
  wire [34:0] _GEN_18 = {{19'd0}, io_data_main_20}; // @[CNN_POOL.scala 26:32]
  wire [35:0] _T_19 = _T_18 + _GEN_18; // @[CNN_POOL.scala 26:32]
  wire [35:0] _GEN_19 = {{20'd0}, io_data_main_21}; // @[CNN_POOL.scala 26:32]
  wire [36:0] _T_20 = _T_19 + _GEN_19; // @[CNN_POOL.scala 26:32]
  wire [36:0] _GEN_20 = {{21'd0}, io_data_main_22}; // @[CNN_POOL.scala 26:32]
  wire [37:0] _T_21 = _T_20 + _GEN_20; // @[CNN_POOL.scala 26:32]
  wire [37:0] _GEN_21 = {{22'd0}, io_data_main_23}; // @[CNN_POOL.scala 26:32]
  wire [38:0] _T_22 = _T_21 + _GEN_21; // @[CNN_POOL.scala 26:32]
  wire [38:0] _GEN_22 = {{23'd0}, io_data_main_24}; // @[CNN_POOL.scala 26:32]
  wire [39:0] _T_23 = _T_22 + _GEN_22; // @[CNN_POOL.scala 26:32]
  wire [20:0] sum = _T_23[20:0]; // @[CNN_POOL.scala 25:17 26:7]
  wire [18:0] _GEN_23 = {{18'd0}, sum[1]}; // @[CNN_POOL.scala 28:25]
  wire [18:0] div4 = sum[20:2] + _GEN_23; // @[CNN_POOL.scala 28:25]
  wire [41:0] mul_res = sum * 21'h1c71c7; // @[CNN_POOL.scala 31:18]
  wire [41:0] _T_28 = {{24'd0}, mul_res[41:24]}; // @[CNN_POOL.scala 32:23]
  wire [41:0] _GEN_25 = {{41'd0}, mul_res[23]}; // @[CNN_POOL.scala 32:32]
  wire [41:0] div9 = _T_28 + _GEN_25; // @[CNN_POOL.scala 32:32]
  wire [16:0] _GEN_26 = {{16'd0}, sum[3]}; // @[CNN_POOL.scala 34:26]
  wire [16:0] div16 = sum[20:4] + _GEN_26; // @[CNN_POOL.scala 34:26]
  wire [50:0] mul_res1 = sum * 30'h33333333; // @[CNN_POOL.scala 40:19]
  wire [50:0] _T_35 = {{32'd0}, mul_res1[50:32]}; // @[CNN_POOL.scala 41:21]
  wire [50:0] _GEN_28 = {{50'd0}, mul_res1[31]}; // @[CNN_POOL.scala 41:30]
  wire [50:0] _T_38 = _T_35 + _GEN_28; // @[CNN_POOL.scala 41:30]
  wire [18:0] div5 = _T_38[18:0]; // @[CNN_POOL.scala 37:18 41:8]
  wire [48:0] mul_res2 = div5 * 30'h33333333; // @[CNN_POOL.scala 42:20]
  wire [48:0] _T_40 = {{32'd0}, mul_res2[48:32]}; // @[CNN_POOL.scala 43:22]
  wire [48:0] _GEN_30 = {{48'd0}, mul_res2[31]}; // @[CNN_POOL.scala 43:31]
  wire [48:0] _T_43 = _T_40 + _GEN_30; // @[CNN_POOL.scala 43:31]
  wire [16:0] div25 = _T_43[16:0]; // @[CNN_POOL.scala 39:19 43:9]
  wire [15:0] _T_50 = 4'h1 == io_k ? sum[15:0] : 16'h0; // @[Mux.scala 80:57]
  wire [15:0] _T_52 = 4'h2 == io_k ? div4[15:0] : _T_50; // @[Mux.scala 80:57]
  wire [15:0] _T_54 = 4'h3 == io_k ? div9[15:0] : _T_52; // @[Mux.scala 80:57]
  wire [15:0] _T_56 = 4'h4 == io_k ? div16[15:0] : _T_54; // @[Mux.scala 80:57]
  assign io_data_res = 4'h5 == io_k ? div25[15:0] : _T_56; // @[Mux.scala 80:57]
endmodule
module CNNPool(
  input  [3:0]  io_k,
  input  [1:0]  io_agm,
  input  [15:0] io_data_main_0,
  input  [15:0] io_data_main_1,
  input  [15:0] io_data_main_2,
  input  [15:0] io_data_main_3,
  input  [15:0] io_data_main_4,
  input  [15:0] io_data_main_5,
  input  [15:0] io_data_main_6,
  input  [15:0] io_data_main_7,
  input  [15:0] io_data_main_8,
  input  [15:0] io_data_main_9,
  input  [15:0] io_data_main_10,
  input  [15:0] io_data_main_11,
  input  [15:0] io_data_main_12,
  input  [15:0] io_data_main_13,
  input  [15:0] io_data_main_14,
  input  [15:0] io_data_main_15,
  input  [15:0] io_data_main_16,
  input  [15:0] io_data_main_17,
  input  [15:0] io_data_main_18,
  input  [15:0] io_data_main_19,
  input  [15:0] io_data_main_20,
  input  [15:0] io_data_main_21,
  input  [15:0] io_data_main_22,
  input  [15:0] io_data_main_23,
  input  [15:0] io_data_main_24,
  output [63:0] io_pool_res
);
  wire [15:0] pool_max_mdu_io_data_main_0; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_1; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_2; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_3; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_4; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_5; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_6; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_7; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_8; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_9; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_10; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_11; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_12; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_13; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_14; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_15; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_16; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_17; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_18; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_19; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_20; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_21; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_22; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_23; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_main_24; // @[CNN_POOL.scala 70:28]
  wire [15:0] pool_max_mdu_io_data_res; // @[CNN_POOL.scala 70:28]
  wire [3:0] pool_avg_mdu_io_k; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_0; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_1; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_2; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_3; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_4; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_5; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_6; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_7; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_8; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_9; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_10; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_11; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_12; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_13; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_14; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_15; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_16; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_17; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_18; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_19; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_20; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_21; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_22; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_23; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_main_24; // @[CNN_POOL.scala 73:28]
  wire [15:0] pool_avg_mdu_io_data_res; // @[CNN_POOL.scala 73:28]
  wire [15:0] _T_1 = 2'h1 == io_agm ? pool_max_mdu_io_data_res : 16'h0; // @[Mux.scala 80:57]
  wire [15:0] res = 2'h2 == io_agm ? pool_avg_mdu_io_data_res : _T_1; // @[Mux.scala 80:57]
  CNNPoolMax pool_max_mdu ( // @[CNN_POOL.scala 70:28]
    .io_data_main_0(pool_max_mdu_io_data_main_0),
    .io_data_main_1(pool_max_mdu_io_data_main_1),
    .io_data_main_2(pool_max_mdu_io_data_main_2),
    .io_data_main_3(pool_max_mdu_io_data_main_3),
    .io_data_main_4(pool_max_mdu_io_data_main_4),
    .io_data_main_5(pool_max_mdu_io_data_main_5),
    .io_data_main_6(pool_max_mdu_io_data_main_6),
    .io_data_main_7(pool_max_mdu_io_data_main_7),
    .io_data_main_8(pool_max_mdu_io_data_main_8),
    .io_data_main_9(pool_max_mdu_io_data_main_9),
    .io_data_main_10(pool_max_mdu_io_data_main_10),
    .io_data_main_11(pool_max_mdu_io_data_main_11),
    .io_data_main_12(pool_max_mdu_io_data_main_12),
    .io_data_main_13(pool_max_mdu_io_data_main_13),
    .io_data_main_14(pool_max_mdu_io_data_main_14),
    .io_data_main_15(pool_max_mdu_io_data_main_15),
    .io_data_main_16(pool_max_mdu_io_data_main_16),
    .io_data_main_17(pool_max_mdu_io_data_main_17),
    .io_data_main_18(pool_max_mdu_io_data_main_18),
    .io_data_main_19(pool_max_mdu_io_data_main_19),
    .io_data_main_20(pool_max_mdu_io_data_main_20),
    .io_data_main_21(pool_max_mdu_io_data_main_21),
    .io_data_main_22(pool_max_mdu_io_data_main_22),
    .io_data_main_23(pool_max_mdu_io_data_main_23),
    .io_data_main_24(pool_max_mdu_io_data_main_24),
    .io_data_res(pool_max_mdu_io_data_res)
  );
  CNNPoolAvg pool_avg_mdu ( // @[CNN_POOL.scala 73:28]
    .io_k(pool_avg_mdu_io_k),
    .io_data_main_0(pool_avg_mdu_io_data_main_0),
    .io_data_main_1(pool_avg_mdu_io_data_main_1),
    .io_data_main_2(pool_avg_mdu_io_data_main_2),
    .io_data_main_3(pool_avg_mdu_io_data_main_3),
    .io_data_main_4(pool_avg_mdu_io_data_main_4),
    .io_data_main_5(pool_avg_mdu_io_data_main_5),
    .io_data_main_6(pool_avg_mdu_io_data_main_6),
    .io_data_main_7(pool_avg_mdu_io_data_main_7),
    .io_data_main_8(pool_avg_mdu_io_data_main_8),
    .io_data_main_9(pool_avg_mdu_io_data_main_9),
    .io_data_main_10(pool_avg_mdu_io_data_main_10),
    .io_data_main_11(pool_avg_mdu_io_data_main_11),
    .io_data_main_12(pool_avg_mdu_io_data_main_12),
    .io_data_main_13(pool_avg_mdu_io_data_main_13),
    .io_data_main_14(pool_avg_mdu_io_data_main_14),
    .io_data_main_15(pool_avg_mdu_io_data_main_15),
    .io_data_main_16(pool_avg_mdu_io_data_main_16),
    .io_data_main_17(pool_avg_mdu_io_data_main_17),
    .io_data_main_18(pool_avg_mdu_io_data_main_18),
    .io_data_main_19(pool_avg_mdu_io_data_main_19),
    .io_data_main_20(pool_avg_mdu_io_data_main_20),
    .io_data_main_21(pool_avg_mdu_io_data_main_21),
    .io_data_main_22(pool_avg_mdu_io_data_main_22),
    .io_data_main_23(pool_avg_mdu_io_data_main_23),
    .io_data_main_24(pool_avg_mdu_io_data_main_24),
    .io_data_res(pool_avg_mdu_io_data_res)
  );
  assign io_pool_res = {48'h0,res}; // @[Cat.scala 30:58]
  assign pool_max_mdu_io_data_main_0 = io_data_main_0; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_1 = io_data_main_1; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_2 = io_data_main_2; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_3 = io_data_main_3; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_4 = io_data_main_4; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_5 = io_data_main_5; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_6 = io_data_main_6; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_7 = io_data_main_7; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_8 = io_data_main_8; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_9 = io_data_main_9; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_10 = io_data_main_10; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_11 = io_data_main_11; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_12 = io_data_main_12; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_13 = io_data_main_13; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_14 = io_data_main_14; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_15 = io_data_main_15; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_16 = io_data_main_16; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_17 = io_data_main_17; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_18 = io_data_main_18; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_19 = io_data_main_19; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_20 = io_data_main_20; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_21 = io_data_main_21; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_22 = io_data_main_22; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_23 = io_data_main_23; // @[CNN_POOL.scala 71:29]
  assign pool_max_mdu_io_data_main_24 = io_data_main_24; // @[CNN_POOL.scala 71:29]
  assign pool_avg_mdu_io_k = io_k; // @[CNN_POOL.scala 75:21]
  assign pool_avg_mdu_io_data_main_0 = io_data_main_0; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_1 = io_data_main_1; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_2 = io_data_main_2; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_3 = io_data_main_3; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_4 = io_data_main_4; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_5 = io_data_main_5; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_6 = io_data_main_6; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_7 = io_data_main_7; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_8 = io_data_main_8; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_9 = io_data_main_9; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_10 = io_data_main_10; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_11 = io_data_main_11; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_12 = io_data_main_12; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_13 = io_data_main_13; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_14 = io_data_main_14; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_15 = io_data_main_15; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_16 = io_data_main_16; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_17 = io_data_main_17; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_18 = io_data_main_18; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_19 = io_data_main_19; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_20 = io_data_main_20; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_21 = io_data_main_21; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_22 = io_data_main_22; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_23 = io_data_main_23; // @[CNN_POOL.scala 74:29]
  assign pool_avg_mdu_io_data_main_24 = io_data_main_24; // @[CNN_POOL.scala 74:29]
endmodule
module CNNActSub(
  input  [15:0] io_in_data_0,
  input  [15:0] io_in_data_1,
  input  [15:0] io_in_data_2,
  input  [15:0] io_in_data_3,
  input  [15:0] io_in_zero_0,
  input  [15:0] io_in_zero_1,
  input  [15:0] io_in_zero_2,
  input  [15:0] io_in_zero_3,
  output [15:0] io_res_0,
  output [15:0] io_res_1,
  output [15:0] io_res_2,
  output [15:0] io_res_3
);
  assign io_res_0 = io_in_data_0 >= io_in_zero_0 ? io_in_data_0 : io_in_zero_0; // @[CNN_ACT.scala 27:21]
  assign io_res_1 = io_in_data_1 >= io_in_zero_1 ? io_in_data_1 : io_in_zero_1; // @[CNN_ACT.scala 27:21]
  assign io_res_2 = io_in_data_2 >= io_in_zero_2 ? io_in_data_2 : io_in_zero_2; // @[CNN_ACT.scala 27:21]
  assign io_res_3 = io_in_data_3 >= io_in_zero_3 ? io_in_data_3 : io_in_zero_3; // @[CNN_ACT.scala 27:21]
endmodule
module CNNActSub_1(
  input  [7:0] io_in_data_0,
  input  [7:0] io_in_data_1,
  input  [7:0] io_in_data_2,
  input  [7:0] io_in_data_3,
  input  [7:0] io_in_data_4,
  input  [7:0] io_in_data_5,
  input  [7:0] io_in_data_6,
  input  [7:0] io_in_data_7,
  input  [7:0] io_in_zero_0,
  input  [7:0] io_in_zero_1,
  input  [7:0] io_in_zero_2,
  input  [7:0] io_in_zero_3,
  input  [7:0] io_in_zero_4,
  input  [7:0] io_in_zero_5,
  input  [7:0] io_in_zero_6,
  input  [7:0] io_in_zero_7,
  output [7:0] io_res_0,
  output [7:0] io_res_1,
  output [7:0] io_res_2,
  output [7:0] io_res_3,
  output [7:0] io_res_4,
  output [7:0] io_res_5,
  output [7:0] io_res_6,
  output [7:0] io_res_7
);
  assign io_res_0 = io_in_data_0 >= io_in_zero_0 ? io_in_data_0 : io_in_zero_0; // @[CNN_ACT.scala 27:21]
  assign io_res_1 = io_in_data_1 >= io_in_zero_1 ? io_in_data_1 : io_in_zero_1; // @[CNN_ACT.scala 27:21]
  assign io_res_2 = io_in_data_2 >= io_in_zero_2 ? io_in_data_2 : io_in_zero_2; // @[CNN_ACT.scala 27:21]
  assign io_res_3 = io_in_data_3 >= io_in_zero_3 ? io_in_data_3 : io_in_zero_3; // @[CNN_ACT.scala 27:21]
  assign io_res_4 = io_in_data_4 >= io_in_zero_4 ? io_in_data_4 : io_in_zero_4; // @[CNN_ACT.scala 27:21]
  assign io_res_5 = io_in_data_5 >= io_in_zero_5 ? io_in_data_5 : io_in_zero_5; // @[CNN_ACT.scala 27:21]
  assign io_res_6 = io_in_data_6 >= io_in_zero_6 ? io_in_data_6 : io_in_zero_6; // @[CNN_ACT.scala 27:21]
  assign io_res_7 = io_in_data_7 >= io_in_zero_7 ? io_in_data_7 : io_in_zero_7; // @[CNN_ACT.scala 27:21]
endmodule
module CNNActSub_2(
  input  [3:0] io_in_data_0,
  input  [3:0] io_in_data_1,
  input  [3:0] io_in_data_2,
  input  [3:0] io_in_data_3,
  input  [3:0] io_in_data_4,
  input  [3:0] io_in_data_5,
  input  [3:0] io_in_data_6,
  input  [3:0] io_in_data_7,
  input  [3:0] io_in_data_8,
  input  [3:0] io_in_data_9,
  input  [3:0] io_in_data_10,
  input  [3:0] io_in_data_11,
  input  [3:0] io_in_data_12,
  input  [3:0] io_in_data_13,
  input  [3:0] io_in_data_14,
  input  [3:0] io_in_data_15,
  input  [3:0] io_in_zero_0,
  input  [3:0] io_in_zero_1,
  input  [3:0] io_in_zero_2,
  input  [3:0] io_in_zero_3,
  input  [3:0] io_in_zero_4,
  input  [3:0] io_in_zero_5,
  input  [3:0] io_in_zero_6,
  input  [3:0] io_in_zero_7,
  input  [3:0] io_in_zero_8,
  input  [3:0] io_in_zero_9,
  input  [3:0] io_in_zero_10,
  input  [3:0] io_in_zero_11,
  input  [3:0] io_in_zero_12,
  input  [3:0] io_in_zero_13,
  input  [3:0] io_in_zero_14,
  input  [3:0] io_in_zero_15,
  output [3:0] io_res_0,
  output [3:0] io_res_1,
  output [3:0] io_res_2,
  output [3:0] io_res_3,
  output [3:0] io_res_4,
  output [3:0] io_res_5,
  output [3:0] io_res_6,
  output [3:0] io_res_7,
  output [3:0] io_res_8,
  output [3:0] io_res_9,
  output [3:0] io_res_10,
  output [3:0] io_res_11,
  output [3:0] io_res_12,
  output [3:0] io_res_13,
  output [3:0] io_res_14,
  output [3:0] io_res_15
);
  assign io_res_0 = io_in_data_0 >= io_in_zero_0 ? io_in_data_0 : io_in_zero_0; // @[CNN_ACT.scala 27:21]
  assign io_res_1 = io_in_data_1 >= io_in_zero_1 ? io_in_data_1 : io_in_zero_1; // @[CNN_ACT.scala 27:21]
  assign io_res_2 = io_in_data_2 >= io_in_zero_2 ? io_in_data_2 : io_in_zero_2; // @[CNN_ACT.scala 27:21]
  assign io_res_3 = io_in_data_3 >= io_in_zero_3 ? io_in_data_3 : io_in_zero_3; // @[CNN_ACT.scala 27:21]
  assign io_res_4 = io_in_data_4 >= io_in_zero_4 ? io_in_data_4 : io_in_zero_4; // @[CNN_ACT.scala 27:21]
  assign io_res_5 = io_in_data_5 >= io_in_zero_5 ? io_in_data_5 : io_in_zero_5; // @[CNN_ACT.scala 27:21]
  assign io_res_6 = io_in_data_6 >= io_in_zero_6 ? io_in_data_6 : io_in_zero_6; // @[CNN_ACT.scala 27:21]
  assign io_res_7 = io_in_data_7 >= io_in_zero_7 ? io_in_data_7 : io_in_zero_7; // @[CNN_ACT.scala 27:21]
  assign io_res_8 = io_in_data_8 >= io_in_zero_8 ? io_in_data_8 : io_in_zero_8; // @[CNN_ACT.scala 27:21]
  assign io_res_9 = io_in_data_9 >= io_in_zero_9 ? io_in_data_9 : io_in_zero_9; // @[CNN_ACT.scala 27:21]
  assign io_res_10 = io_in_data_10 >= io_in_zero_10 ? io_in_data_10 : io_in_zero_10; // @[CNN_ACT.scala 27:21]
  assign io_res_11 = io_in_data_11 >= io_in_zero_11 ? io_in_data_11 : io_in_zero_11; // @[CNN_ACT.scala 27:21]
  assign io_res_12 = io_in_data_12 >= io_in_zero_12 ? io_in_data_12 : io_in_zero_12; // @[CNN_ACT.scala 27:21]
  assign io_res_13 = io_in_data_13 >= io_in_zero_13 ? io_in_data_13 : io_in_zero_13; // @[CNN_ACT.scala 27:21]
  assign io_res_14 = io_in_data_14 >= io_in_zero_14 ? io_in_data_14 : io_in_zero_14; // @[CNN_ACT.scala 27:21]
  assign io_res_15 = io_in_data_15 >= io_in_zero_15 ? io_in_data_15 : io_in_zero_15; // @[CNN_ACT.scala 27:21]
endmodule
module CNNActSub_3(
  input  [1:0] io_in_data_0,
  input  [1:0] io_in_data_1,
  input  [1:0] io_in_data_2,
  input  [1:0] io_in_data_3,
  input  [1:0] io_in_data_4,
  input  [1:0] io_in_data_5,
  input  [1:0] io_in_data_6,
  input  [1:0] io_in_data_7,
  input  [1:0] io_in_data_8,
  input  [1:0] io_in_data_9,
  input  [1:0] io_in_data_10,
  input  [1:0] io_in_data_11,
  input  [1:0] io_in_data_12,
  input  [1:0] io_in_data_13,
  input  [1:0] io_in_data_14,
  input  [1:0] io_in_data_15,
  input  [1:0] io_in_data_16,
  input  [1:0] io_in_data_17,
  input  [1:0] io_in_data_18,
  input  [1:0] io_in_data_19,
  input  [1:0] io_in_data_20,
  input  [1:0] io_in_data_21,
  input  [1:0] io_in_data_22,
  input  [1:0] io_in_data_23,
  input  [1:0] io_in_data_24,
  input  [1:0] io_in_data_25,
  input  [1:0] io_in_data_26,
  input  [1:0] io_in_data_27,
  input  [1:0] io_in_data_28,
  input  [1:0] io_in_data_29,
  input  [1:0] io_in_data_30,
  input  [1:0] io_in_data_31,
  input  [1:0] io_in_zero_0,
  input  [1:0] io_in_zero_1,
  input  [1:0] io_in_zero_2,
  input  [1:0] io_in_zero_3,
  input  [1:0] io_in_zero_4,
  input  [1:0] io_in_zero_5,
  input  [1:0] io_in_zero_6,
  input  [1:0] io_in_zero_7,
  input  [1:0] io_in_zero_8,
  input  [1:0] io_in_zero_9,
  input  [1:0] io_in_zero_10,
  input  [1:0] io_in_zero_11,
  input  [1:0] io_in_zero_12,
  input  [1:0] io_in_zero_13,
  input  [1:0] io_in_zero_14,
  input  [1:0] io_in_zero_15,
  input  [1:0] io_in_zero_16,
  input  [1:0] io_in_zero_17,
  input  [1:0] io_in_zero_18,
  input  [1:0] io_in_zero_19,
  input  [1:0] io_in_zero_20,
  input  [1:0] io_in_zero_21,
  input  [1:0] io_in_zero_22,
  input  [1:0] io_in_zero_23,
  input  [1:0] io_in_zero_24,
  input  [1:0] io_in_zero_25,
  input  [1:0] io_in_zero_26,
  input  [1:0] io_in_zero_27,
  input  [1:0] io_in_zero_28,
  input  [1:0] io_in_zero_29,
  input  [1:0] io_in_zero_30,
  input  [1:0] io_in_zero_31,
  output [1:0] io_res_0,
  output [1:0] io_res_1,
  output [1:0] io_res_2,
  output [1:0] io_res_3,
  output [1:0] io_res_4,
  output [1:0] io_res_5,
  output [1:0] io_res_6,
  output [1:0] io_res_7,
  output [1:0] io_res_8,
  output [1:0] io_res_9,
  output [1:0] io_res_10,
  output [1:0] io_res_11,
  output [1:0] io_res_12,
  output [1:0] io_res_13,
  output [1:0] io_res_14,
  output [1:0] io_res_15,
  output [1:0] io_res_16,
  output [1:0] io_res_17,
  output [1:0] io_res_18,
  output [1:0] io_res_19,
  output [1:0] io_res_20,
  output [1:0] io_res_21,
  output [1:0] io_res_22,
  output [1:0] io_res_23,
  output [1:0] io_res_24,
  output [1:0] io_res_25,
  output [1:0] io_res_26,
  output [1:0] io_res_27,
  output [1:0] io_res_28,
  output [1:0] io_res_29,
  output [1:0] io_res_30,
  output [1:0] io_res_31
);
  assign io_res_0 = io_in_data_0 >= io_in_zero_0 ? io_in_data_0 : io_in_zero_0; // @[CNN_ACT.scala 27:21]
  assign io_res_1 = io_in_data_1 >= io_in_zero_1 ? io_in_data_1 : io_in_zero_1; // @[CNN_ACT.scala 27:21]
  assign io_res_2 = io_in_data_2 >= io_in_zero_2 ? io_in_data_2 : io_in_zero_2; // @[CNN_ACT.scala 27:21]
  assign io_res_3 = io_in_data_3 >= io_in_zero_3 ? io_in_data_3 : io_in_zero_3; // @[CNN_ACT.scala 27:21]
  assign io_res_4 = io_in_data_4 >= io_in_zero_4 ? io_in_data_4 : io_in_zero_4; // @[CNN_ACT.scala 27:21]
  assign io_res_5 = io_in_data_5 >= io_in_zero_5 ? io_in_data_5 : io_in_zero_5; // @[CNN_ACT.scala 27:21]
  assign io_res_6 = io_in_data_6 >= io_in_zero_6 ? io_in_data_6 : io_in_zero_6; // @[CNN_ACT.scala 27:21]
  assign io_res_7 = io_in_data_7 >= io_in_zero_7 ? io_in_data_7 : io_in_zero_7; // @[CNN_ACT.scala 27:21]
  assign io_res_8 = io_in_data_8 >= io_in_zero_8 ? io_in_data_8 : io_in_zero_8; // @[CNN_ACT.scala 27:21]
  assign io_res_9 = io_in_data_9 >= io_in_zero_9 ? io_in_data_9 : io_in_zero_9; // @[CNN_ACT.scala 27:21]
  assign io_res_10 = io_in_data_10 >= io_in_zero_10 ? io_in_data_10 : io_in_zero_10; // @[CNN_ACT.scala 27:21]
  assign io_res_11 = io_in_data_11 >= io_in_zero_11 ? io_in_data_11 : io_in_zero_11; // @[CNN_ACT.scala 27:21]
  assign io_res_12 = io_in_data_12 >= io_in_zero_12 ? io_in_data_12 : io_in_zero_12; // @[CNN_ACT.scala 27:21]
  assign io_res_13 = io_in_data_13 >= io_in_zero_13 ? io_in_data_13 : io_in_zero_13; // @[CNN_ACT.scala 27:21]
  assign io_res_14 = io_in_data_14 >= io_in_zero_14 ? io_in_data_14 : io_in_zero_14; // @[CNN_ACT.scala 27:21]
  assign io_res_15 = io_in_data_15 >= io_in_zero_15 ? io_in_data_15 : io_in_zero_15; // @[CNN_ACT.scala 27:21]
  assign io_res_16 = io_in_data_16 >= io_in_zero_16 ? io_in_data_16 : io_in_zero_16; // @[CNN_ACT.scala 27:21]
  assign io_res_17 = io_in_data_17 >= io_in_zero_17 ? io_in_data_17 : io_in_zero_17; // @[CNN_ACT.scala 27:21]
  assign io_res_18 = io_in_data_18 >= io_in_zero_18 ? io_in_data_18 : io_in_zero_18; // @[CNN_ACT.scala 27:21]
  assign io_res_19 = io_in_data_19 >= io_in_zero_19 ? io_in_data_19 : io_in_zero_19; // @[CNN_ACT.scala 27:21]
  assign io_res_20 = io_in_data_20 >= io_in_zero_20 ? io_in_data_20 : io_in_zero_20; // @[CNN_ACT.scala 27:21]
  assign io_res_21 = io_in_data_21 >= io_in_zero_21 ? io_in_data_21 : io_in_zero_21; // @[CNN_ACT.scala 27:21]
  assign io_res_22 = io_in_data_22 >= io_in_zero_22 ? io_in_data_22 : io_in_zero_22; // @[CNN_ACT.scala 27:21]
  assign io_res_23 = io_in_data_23 >= io_in_zero_23 ? io_in_data_23 : io_in_zero_23; // @[CNN_ACT.scala 27:21]
  assign io_res_24 = io_in_data_24 >= io_in_zero_24 ? io_in_data_24 : io_in_zero_24; // @[CNN_ACT.scala 27:21]
  assign io_res_25 = io_in_data_25 >= io_in_zero_25 ? io_in_data_25 : io_in_zero_25; // @[CNN_ACT.scala 27:21]
  assign io_res_26 = io_in_data_26 >= io_in_zero_26 ? io_in_data_26 : io_in_zero_26; // @[CNN_ACT.scala 27:21]
  assign io_res_27 = io_in_data_27 >= io_in_zero_27 ? io_in_data_27 : io_in_zero_27; // @[CNN_ACT.scala 27:21]
  assign io_res_28 = io_in_data_28 >= io_in_zero_28 ? io_in_data_28 : io_in_zero_28; // @[CNN_ACT.scala 27:21]
  assign io_res_29 = io_in_data_29 >= io_in_zero_29 ? io_in_data_29 : io_in_zero_29; // @[CNN_ACT.scala 27:21]
  assign io_res_30 = io_in_data_30 >= io_in_zero_30 ? io_in_data_30 : io_in_zero_30; // @[CNN_ACT.scala 27:21]
  assign io_res_31 = io_in_data_31 >= io_in_zero_31 ? io_in_data_31 : io_in_zero_31; // @[CNN_ACT.scala 27:21]
endmodule
module CNNAct(
  input  [63:0] io_data_main,
  input  [63:0] io_data_zero,
  input  [3:0]  io_data_vwidth,
  output [63:0] io_act_res
);
  wire [15:0] act_mdu_4_16_io_in_data_0; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_in_data_1; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_in_data_2; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_in_data_3; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_in_zero_0; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_in_zero_1; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_in_zero_2; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_in_zero_3; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_res_0; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_res_1; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_res_2; // @[CNN_ACT.scala 34:28]
  wire [15:0] act_mdu_4_16_io_res_3; // @[CNN_ACT.scala 34:28]
  wire [7:0] act_mdu_8_8_io_in_data_0; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_data_1; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_data_2; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_data_3; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_data_4; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_data_5; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_data_6; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_data_7; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_0; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_1; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_2; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_3; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_4; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_5; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_6; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_in_zero_7; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_0; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_1; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_2; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_3; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_4; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_5; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_6; // @[CNN_ACT.scala 40:27]
  wire [7:0] act_mdu_8_8_io_res_7; // @[CNN_ACT.scala 40:27]
  wire [3:0] act_mdu_16_4_io_in_data_0; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_1; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_2; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_3; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_4; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_5; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_6; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_7; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_8; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_9; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_10; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_11; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_12; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_13; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_14; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_data_15; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_0; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_1; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_2; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_3; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_4; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_5; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_6; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_7; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_8; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_9; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_10; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_11; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_12; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_13; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_14; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_in_zero_15; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_0; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_1; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_2; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_3; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_4; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_5; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_6; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_7; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_8; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_9; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_10; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_11; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_12; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_13; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_14; // @[CNN_ACT.scala 46:28]
  wire [3:0] act_mdu_16_4_io_res_15; // @[CNN_ACT.scala 46:28]
  wire [1:0] act_mdu_32_2_io_in_data_0; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_1; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_2; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_3; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_4; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_5; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_6; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_7; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_8; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_9; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_10; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_11; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_12; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_13; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_14; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_15; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_16; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_17; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_18; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_19; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_20; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_21; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_22; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_23; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_24; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_25; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_26; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_27; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_28; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_29; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_30; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_data_31; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_0; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_1; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_2; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_3; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_4; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_5; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_6; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_7; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_8; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_9; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_10; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_11; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_12; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_13; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_14; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_15; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_16; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_17; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_18; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_19; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_20; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_21; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_22; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_23; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_24; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_25; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_26; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_27; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_28; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_29; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_30; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_in_zero_31; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_0; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_1; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_2; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_3; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_4; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_5; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_6; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_7; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_8; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_9; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_10; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_11; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_12; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_13; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_14; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_15; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_16; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_17; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_18; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_19; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_20; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_21; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_22; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_23; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_24; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_25; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_26; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_27; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_28; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_29; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_30; // @[CNN_ACT.scala 52:28]
  wire [1:0] act_mdu_32_2_io_res_31; // @[CNN_ACT.scala 52:28]
  wire [63:0] _T_122 = {act_mdu_4_16_io_res_3,act_mdu_4_16_io_res_2,act_mdu_4_16_io_res_1,act_mdu_4_16_io_res_0}; // @[Cat.scala 30:58]
  wire [63:0] _T_129 = {act_mdu_8_8_io_res_7,act_mdu_8_8_io_res_6,act_mdu_8_8_io_res_5,act_mdu_8_8_io_res_4,
    act_mdu_8_8_io_res_3,act_mdu_8_8_io_res_2,act_mdu_8_8_io_res_1,act_mdu_8_8_io_res_0}; // @[Cat.scala 30:58]
  wire [39:0] _T_138 = {act_mdu_16_4_io_res_9,act_mdu_16_4_io_res_8,act_mdu_16_4_io_res_7,act_mdu_16_4_io_res_6,
    act_mdu_16_4_io_res_5,act_mdu_16_4_io_res_4,act_mdu_16_4_io_res_3,act_mdu_16_4_io_res_2,act_mdu_16_4_io_res_1,
    act_mdu_16_4_io_res_0}; // @[Cat.scala 30:58]
  wire [63:0] _T_144 = {act_mdu_16_4_io_res_15,act_mdu_16_4_io_res_14,act_mdu_16_4_io_res_13,act_mdu_16_4_io_res_12,
    act_mdu_16_4_io_res_11,act_mdu_16_4_io_res_10,_T_138}; // @[Cat.scala 30:58]
  wire [19:0] _T_153 = {act_mdu_32_2_io_res_9,act_mdu_32_2_io_res_8,act_mdu_32_2_io_res_7,act_mdu_32_2_io_res_6,
    act_mdu_32_2_io_res_5,act_mdu_32_2_io_res_4,act_mdu_32_2_io_res_3,act_mdu_32_2_io_res_2,act_mdu_32_2_io_res_1,
    act_mdu_32_2_io_res_0}; // @[Cat.scala 30:58]
  wire [37:0] _T_162 = {act_mdu_32_2_io_res_18,act_mdu_32_2_io_res_17,act_mdu_32_2_io_res_16,act_mdu_32_2_io_res_15,
    act_mdu_32_2_io_res_14,act_mdu_32_2_io_res_13,act_mdu_32_2_io_res_12,act_mdu_32_2_io_res_11,act_mdu_32_2_io_res_10,
    _T_153}; // @[Cat.scala 30:58]
  wire [55:0] _T_171 = {act_mdu_32_2_io_res_27,act_mdu_32_2_io_res_26,act_mdu_32_2_io_res_25,act_mdu_32_2_io_res_24,
    act_mdu_32_2_io_res_23,act_mdu_32_2_io_res_22,act_mdu_32_2_io_res_21,act_mdu_32_2_io_res_20,act_mdu_32_2_io_res_19,
    _T_162}; // @[Cat.scala 30:58]
  wire [63:0] _T_175 = {act_mdu_32_2_io_res_31,act_mdu_32_2_io_res_30,act_mdu_32_2_io_res_29,act_mdu_32_2_io_res_28,
    _T_171}; // @[Cat.scala 30:58]
  wire [63:0] _T_177 = 4'h8 == io_data_vwidth ? _T_122 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_179 = 4'h4 == io_data_vwidth ? _T_129 : _T_177; // @[Mux.scala 80:57]
  wire [63:0] _T_181 = 4'h2 == io_data_vwidth ? _T_144 : _T_179; // @[Mux.scala 80:57]
  CNNActSub act_mdu_4_16 ( // @[CNN_ACT.scala 34:28]
    .io_in_data_0(act_mdu_4_16_io_in_data_0),
    .io_in_data_1(act_mdu_4_16_io_in_data_1),
    .io_in_data_2(act_mdu_4_16_io_in_data_2),
    .io_in_data_3(act_mdu_4_16_io_in_data_3),
    .io_in_zero_0(act_mdu_4_16_io_in_zero_0),
    .io_in_zero_1(act_mdu_4_16_io_in_zero_1),
    .io_in_zero_2(act_mdu_4_16_io_in_zero_2),
    .io_in_zero_3(act_mdu_4_16_io_in_zero_3),
    .io_res_0(act_mdu_4_16_io_res_0),
    .io_res_1(act_mdu_4_16_io_res_1),
    .io_res_2(act_mdu_4_16_io_res_2),
    .io_res_3(act_mdu_4_16_io_res_3)
  );
  CNNActSub_1 act_mdu_8_8 ( // @[CNN_ACT.scala 40:27]
    .io_in_data_0(act_mdu_8_8_io_in_data_0),
    .io_in_data_1(act_mdu_8_8_io_in_data_1),
    .io_in_data_2(act_mdu_8_8_io_in_data_2),
    .io_in_data_3(act_mdu_8_8_io_in_data_3),
    .io_in_data_4(act_mdu_8_8_io_in_data_4),
    .io_in_data_5(act_mdu_8_8_io_in_data_5),
    .io_in_data_6(act_mdu_8_8_io_in_data_6),
    .io_in_data_7(act_mdu_8_8_io_in_data_7),
    .io_in_zero_0(act_mdu_8_8_io_in_zero_0),
    .io_in_zero_1(act_mdu_8_8_io_in_zero_1),
    .io_in_zero_2(act_mdu_8_8_io_in_zero_2),
    .io_in_zero_3(act_mdu_8_8_io_in_zero_3),
    .io_in_zero_4(act_mdu_8_8_io_in_zero_4),
    .io_in_zero_5(act_mdu_8_8_io_in_zero_5),
    .io_in_zero_6(act_mdu_8_8_io_in_zero_6),
    .io_in_zero_7(act_mdu_8_8_io_in_zero_7),
    .io_res_0(act_mdu_8_8_io_res_0),
    .io_res_1(act_mdu_8_8_io_res_1),
    .io_res_2(act_mdu_8_8_io_res_2),
    .io_res_3(act_mdu_8_8_io_res_3),
    .io_res_4(act_mdu_8_8_io_res_4),
    .io_res_5(act_mdu_8_8_io_res_5),
    .io_res_6(act_mdu_8_8_io_res_6),
    .io_res_7(act_mdu_8_8_io_res_7)
  );
  CNNActSub_2 act_mdu_16_4 ( // @[CNN_ACT.scala 46:28]
    .io_in_data_0(act_mdu_16_4_io_in_data_0),
    .io_in_data_1(act_mdu_16_4_io_in_data_1),
    .io_in_data_2(act_mdu_16_4_io_in_data_2),
    .io_in_data_3(act_mdu_16_4_io_in_data_3),
    .io_in_data_4(act_mdu_16_4_io_in_data_4),
    .io_in_data_5(act_mdu_16_4_io_in_data_5),
    .io_in_data_6(act_mdu_16_4_io_in_data_6),
    .io_in_data_7(act_mdu_16_4_io_in_data_7),
    .io_in_data_8(act_mdu_16_4_io_in_data_8),
    .io_in_data_9(act_mdu_16_4_io_in_data_9),
    .io_in_data_10(act_mdu_16_4_io_in_data_10),
    .io_in_data_11(act_mdu_16_4_io_in_data_11),
    .io_in_data_12(act_mdu_16_4_io_in_data_12),
    .io_in_data_13(act_mdu_16_4_io_in_data_13),
    .io_in_data_14(act_mdu_16_4_io_in_data_14),
    .io_in_data_15(act_mdu_16_4_io_in_data_15),
    .io_in_zero_0(act_mdu_16_4_io_in_zero_0),
    .io_in_zero_1(act_mdu_16_4_io_in_zero_1),
    .io_in_zero_2(act_mdu_16_4_io_in_zero_2),
    .io_in_zero_3(act_mdu_16_4_io_in_zero_3),
    .io_in_zero_4(act_mdu_16_4_io_in_zero_4),
    .io_in_zero_5(act_mdu_16_4_io_in_zero_5),
    .io_in_zero_6(act_mdu_16_4_io_in_zero_6),
    .io_in_zero_7(act_mdu_16_4_io_in_zero_7),
    .io_in_zero_8(act_mdu_16_4_io_in_zero_8),
    .io_in_zero_9(act_mdu_16_4_io_in_zero_9),
    .io_in_zero_10(act_mdu_16_4_io_in_zero_10),
    .io_in_zero_11(act_mdu_16_4_io_in_zero_11),
    .io_in_zero_12(act_mdu_16_4_io_in_zero_12),
    .io_in_zero_13(act_mdu_16_4_io_in_zero_13),
    .io_in_zero_14(act_mdu_16_4_io_in_zero_14),
    .io_in_zero_15(act_mdu_16_4_io_in_zero_15),
    .io_res_0(act_mdu_16_4_io_res_0),
    .io_res_1(act_mdu_16_4_io_res_1),
    .io_res_2(act_mdu_16_4_io_res_2),
    .io_res_3(act_mdu_16_4_io_res_3),
    .io_res_4(act_mdu_16_4_io_res_4),
    .io_res_5(act_mdu_16_4_io_res_5),
    .io_res_6(act_mdu_16_4_io_res_6),
    .io_res_7(act_mdu_16_4_io_res_7),
    .io_res_8(act_mdu_16_4_io_res_8),
    .io_res_9(act_mdu_16_4_io_res_9),
    .io_res_10(act_mdu_16_4_io_res_10),
    .io_res_11(act_mdu_16_4_io_res_11),
    .io_res_12(act_mdu_16_4_io_res_12),
    .io_res_13(act_mdu_16_4_io_res_13),
    .io_res_14(act_mdu_16_4_io_res_14),
    .io_res_15(act_mdu_16_4_io_res_15)
  );
  CNNActSub_3 act_mdu_32_2 ( // @[CNN_ACT.scala 52:28]
    .io_in_data_0(act_mdu_32_2_io_in_data_0),
    .io_in_data_1(act_mdu_32_2_io_in_data_1),
    .io_in_data_2(act_mdu_32_2_io_in_data_2),
    .io_in_data_3(act_mdu_32_2_io_in_data_3),
    .io_in_data_4(act_mdu_32_2_io_in_data_4),
    .io_in_data_5(act_mdu_32_2_io_in_data_5),
    .io_in_data_6(act_mdu_32_2_io_in_data_6),
    .io_in_data_7(act_mdu_32_2_io_in_data_7),
    .io_in_data_8(act_mdu_32_2_io_in_data_8),
    .io_in_data_9(act_mdu_32_2_io_in_data_9),
    .io_in_data_10(act_mdu_32_2_io_in_data_10),
    .io_in_data_11(act_mdu_32_2_io_in_data_11),
    .io_in_data_12(act_mdu_32_2_io_in_data_12),
    .io_in_data_13(act_mdu_32_2_io_in_data_13),
    .io_in_data_14(act_mdu_32_2_io_in_data_14),
    .io_in_data_15(act_mdu_32_2_io_in_data_15),
    .io_in_data_16(act_mdu_32_2_io_in_data_16),
    .io_in_data_17(act_mdu_32_2_io_in_data_17),
    .io_in_data_18(act_mdu_32_2_io_in_data_18),
    .io_in_data_19(act_mdu_32_2_io_in_data_19),
    .io_in_data_20(act_mdu_32_2_io_in_data_20),
    .io_in_data_21(act_mdu_32_2_io_in_data_21),
    .io_in_data_22(act_mdu_32_2_io_in_data_22),
    .io_in_data_23(act_mdu_32_2_io_in_data_23),
    .io_in_data_24(act_mdu_32_2_io_in_data_24),
    .io_in_data_25(act_mdu_32_2_io_in_data_25),
    .io_in_data_26(act_mdu_32_2_io_in_data_26),
    .io_in_data_27(act_mdu_32_2_io_in_data_27),
    .io_in_data_28(act_mdu_32_2_io_in_data_28),
    .io_in_data_29(act_mdu_32_2_io_in_data_29),
    .io_in_data_30(act_mdu_32_2_io_in_data_30),
    .io_in_data_31(act_mdu_32_2_io_in_data_31),
    .io_in_zero_0(act_mdu_32_2_io_in_zero_0),
    .io_in_zero_1(act_mdu_32_2_io_in_zero_1),
    .io_in_zero_2(act_mdu_32_2_io_in_zero_2),
    .io_in_zero_3(act_mdu_32_2_io_in_zero_3),
    .io_in_zero_4(act_mdu_32_2_io_in_zero_4),
    .io_in_zero_5(act_mdu_32_2_io_in_zero_5),
    .io_in_zero_6(act_mdu_32_2_io_in_zero_6),
    .io_in_zero_7(act_mdu_32_2_io_in_zero_7),
    .io_in_zero_8(act_mdu_32_2_io_in_zero_8),
    .io_in_zero_9(act_mdu_32_2_io_in_zero_9),
    .io_in_zero_10(act_mdu_32_2_io_in_zero_10),
    .io_in_zero_11(act_mdu_32_2_io_in_zero_11),
    .io_in_zero_12(act_mdu_32_2_io_in_zero_12),
    .io_in_zero_13(act_mdu_32_2_io_in_zero_13),
    .io_in_zero_14(act_mdu_32_2_io_in_zero_14),
    .io_in_zero_15(act_mdu_32_2_io_in_zero_15),
    .io_in_zero_16(act_mdu_32_2_io_in_zero_16),
    .io_in_zero_17(act_mdu_32_2_io_in_zero_17),
    .io_in_zero_18(act_mdu_32_2_io_in_zero_18),
    .io_in_zero_19(act_mdu_32_2_io_in_zero_19),
    .io_in_zero_20(act_mdu_32_2_io_in_zero_20),
    .io_in_zero_21(act_mdu_32_2_io_in_zero_21),
    .io_in_zero_22(act_mdu_32_2_io_in_zero_22),
    .io_in_zero_23(act_mdu_32_2_io_in_zero_23),
    .io_in_zero_24(act_mdu_32_2_io_in_zero_24),
    .io_in_zero_25(act_mdu_32_2_io_in_zero_25),
    .io_in_zero_26(act_mdu_32_2_io_in_zero_26),
    .io_in_zero_27(act_mdu_32_2_io_in_zero_27),
    .io_in_zero_28(act_mdu_32_2_io_in_zero_28),
    .io_in_zero_29(act_mdu_32_2_io_in_zero_29),
    .io_in_zero_30(act_mdu_32_2_io_in_zero_30),
    .io_in_zero_31(act_mdu_32_2_io_in_zero_31),
    .io_res_0(act_mdu_32_2_io_res_0),
    .io_res_1(act_mdu_32_2_io_res_1),
    .io_res_2(act_mdu_32_2_io_res_2),
    .io_res_3(act_mdu_32_2_io_res_3),
    .io_res_4(act_mdu_32_2_io_res_4),
    .io_res_5(act_mdu_32_2_io_res_5),
    .io_res_6(act_mdu_32_2_io_res_6),
    .io_res_7(act_mdu_32_2_io_res_7),
    .io_res_8(act_mdu_32_2_io_res_8),
    .io_res_9(act_mdu_32_2_io_res_9),
    .io_res_10(act_mdu_32_2_io_res_10),
    .io_res_11(act_mdu_32_2_io_res_11),
    .io_res_12(act_mdu_32_2_io_res_12),
    .io_res_13(act_mdu_32_2_io_res_13),
    .io_res_14(act_mdu_32_2_io_res_14),
    .io_res_15(act_mdu_32_2_io_res_15),
    .io_res_16(act_mdu_32_2_io_res_16),
    .io_res_17(act_mdu_32_2_io_res_17),
    .io_res_18(act_mdu_32_2_io_res_18),
    .io_res_19(act_mdu_32_2_io_res_19),
    .io_res_20(act_mdu_32_2_io_res_20),
    .io_res_21(act_mdu_32_2_io_res_21),
    .io_res_22(act_mdu_32_2_io_res_22),
    .io_res_23(act_mdu_32_2_io_res_23),
    .io_res_24(act_mdu_32_2_io_res_24),
    .io_res_25(act_mdu_32_2_io_res_25),
    .io_res_26(act_mdu_32_2_io_res_26),
    .io_res_27(act_mdu_32_2_io_res_27),
    .io_res_28(act_mdu_32_2_io_res_28),
    .io_res_29(act_mdu_32_2_io_res_29),
    .io_res_30(act_mdu_32_2_io_res_30),
    .io_res_31(act_mdu_32_2_io_res_31)
  );
  assign io_act_res = 4'h1 == io_data_vwidth ? _T_175 : _T_181; // @[Mux.scala 80:57]
  assign act_mdu_4_16_io_in_data_0 = io_data_main[15:0]; // @[CNN_ACT.scala 36:47]
  assign act_mdu_4_16_io_in_data_1 = io_data_main[31:16]; // @[CNN_ACT.scala 36:47]
  assign act_mdu_4_16_io_in_data_2 = io_data_main[47:32]; // @[CNN_ACT.scala 36:47]
  assign act_mdu_4_16_io_in_data_3 = io_data_main[63:48]; // @[CNN_ACT.scala 36:47]
  assign act_mdu_4_16_io_in_zero_0 = io_data_zero[15:0]; // @[CNN_ACT.scala 37:47]
  assign act_mdu_4_16_io_in_zero_1 = io_data_zero[31:16]; // @[CNN_ACT.scala 37:47]
  assign act_mdu_4_16_io_in_zero_2 = io_data_zero[47:32]; // @[CNN_ACT.scala 37:47]
  assign act_mdu_4_16_io_in_zero_3 = io_data_zero[63:48]; // @[CNN_ACT.scala 37:47]
  assign act_mdu_8_8_io_in_data_0 = io_data_main[7:0]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_data_1 = io_data_main[15:8]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_data_2 = io_data_main[23:16]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_data_3 = io_data_main[31:24]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_data_4 = io_data_main[39:32]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_data_5 = io_data_main[47:40]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_data_6 = io_data_main[55:48]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_data_7 = io_data_main[63:56]; // @[CNN_ACT.scala 42:46]
  assign act_mdu_8_8_io_in_zero_0 = io_data_zero[7:0]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_8_8_io_in_zero_1 = io_data_zero[15:8]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_8_8_io_in_zero_2 = io_data_zero[23:16]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_8_8_io_in_zero_3 = io_data_zero[31:24]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_8_8_io_in_zero_4 = io_data_zero[39:32]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_8_8_io_in_zero_5 = io_data_zero[47:40]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_8_8_io_in_zero_6 = io_data_zero[55:48]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_8_8_io_in_zero_7 = io_data_zero[63:56]; // @[CNN_ACT.scala 43:46]
  assign act_mdu_16_4_io_in_data_0 = io_data_main[3:0]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_1 = io_data_main[7:4]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_2 = io_data_main[11:8]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_3 = io_data_main[15:12]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_4 = io_data_main[19:16]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_5 = io_data_main[23:20]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_6 = io_data_main[27:24]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_7 = io_data_main[31:28]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_8 = io_data_main[35:32]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_9 = io_data_main[39:36]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_10 = io_data_main[43:40]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_11 = io_data_main[47:44]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_12 = io_data_main[51:48]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_13 = io_data_main[55:52]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_14 = io_data_main[59:56]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_data_15 = io_data_main[63:60]; // @[CNN_ACT.scala 48:47]
  assign act_mdu_16_4_io_in_zero_0 = io_data_zero[3:0]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_1 = io_data_zero[7:4]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_2 = io_data_zero[11:8]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_3 = io_data_zero[15:12]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_4 = io_data_zero[19:16]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_5 = io_data_zero[23:20]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_6 = io_data_zero[27:24]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_7 = io_data_zero[31:28]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_8 = io_data_zero[35:32]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_9 = io_data_zero[39:36]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_10 = io_data_zero[43:40]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_11 = io_data_zero[47:44]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_12 = io_data_zero[51:48]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_13 = io_data_zero[55:52]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_14 = io_data_zero[59:56]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_16_4_io_in_zero_15 = io_data_zero[63:60]; // @[CNN_ACT.scala 49:47]
  assign act_mdu_32_2_io_in_data_0 = io_data_main[1:0]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_1 = io_data_main[3:2]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_2 = io_data_main[5:4]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_3 = io_data_main[7:6]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_4 = io_data_main[9:8]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_5 = io_data_main[11:10]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_6 = io_data_main[13:12]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_7 = io_data_main[15:14]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_8 = io_data_main[17:16]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_9 = io_data_main[19:18]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_10 = io_data_main[21:20]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_11 = io_data_main[23:22]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_12 = io_data_main[25:24]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_13 = io_data_main[27:26]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_14 = io_data_main[29:28]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_15 = io_data_main[31:30]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_16 = io_data_main[33:32]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_17 = io_data_main[35:34]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_18 = io_data_main[37:36]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_19 = io_data_main[39:38]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_20 = io_data_main[41:40]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_21 = io_data_main[43:42]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_22 = io_data_main[45:44]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_23 = io_data_main[47:46]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_24 = io_data_main[49:48]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_25 = io_data_main[51:50]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_26 = io_data_main[53:52]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_27 = io_data_main[55:54]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_28 = io_data_main[57:56]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_29 = io_data_main[59:58]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_30 = io_data_main[61:60]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_data_31 = io_data_main[63:62]; // @[CNN_ACT.scala 54:47]
  assign act_mdu_32_2_io_in_zero_0 = io_data_zero[1:0]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_1 = io_data_zero[3:2]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_2 = io_data_zero[5:4]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_3 = io_data_zero[7:6]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_4 = io_data_zero[9:8]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_5 = io_data_zero[11:10]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_6 = io_data_zero[13:12]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_7 = io_data_zero[15:14]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_8 = io_data_zero[17:16]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_9 = io_data_zero[19:18]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_10 = io_data_zero[21:20]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_11 = io_data_zero[23:22]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_12 = io_data_zero[25:24]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_13 = io_data_zero[27:26]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_14 = io_data_zero[29:28]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_15 = io_data_zero[31:30]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_16 = io_data_zero[33:32]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_17 = io_data_zero[35:34]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_18 = io_data_zero[37:36]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_19 = io_data_zero[39:38]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_20 = io_data_zero[41:40]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_21 = io_data_zero[43:42]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_22 = io_data_zero[45:44]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_23 = io_data_zero[47:46]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_24 = io_data_zero[49:48]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_25 = io_data_zero[51:50]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_26 = io_data_zero[53:52]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_27 = io_data_zero[55:54]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_28 = io_data_zero[57:56]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_29 = io_data_zero[59:58]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_30 = io_data_zero[61:60]; // @[CNN_ACT.scala 55:47]
  assign act_mdu_32_2_io_in_zero_31 = io_data_zero[63:62]; // @[CNN_ACT.scala 55:47]
endmodule
module CNNFU(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_imm,
  input  [2:0]  io_vtag,
  input  [3:0]  io_length_k,
  input  [4:0]  io_vec_addr,
  input  [1:0]  io_algorithm,
  output        io_loadv_valid,
  output [63:0] io_loadv_src1,
  output [63:0] io_loadv_src2,
  output [6:0]  io_loadv_func,
  input         io_loadv_load_valid,
  input  [63:0] io_loadv_load_data,
  input         io_loadv_load_exception
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  vreg_mdu_clock; // @[CNN_FU.scala 86:24]
  wire [4:0] vreg_mdu_io_vaddr; // @[CNN_FU.scala 86:24]
  wire [2:0] vreg_mdu_io_vtag; // @[CNN_FU.scala 86:24]
  wire [2:0] vreg_mdu_io_vop; // @[CNN_FU.scala 86:24]
  wire [3:0] vreg_mdu_io_k; // @[CNN_FU.scala 86:24]
  wire  vreg_mdu_io_vwen; // @[CNN_FU.scala 86:24]
  wire [79:0] vreg_mdu_io_load_data; // @[CNN_FU.scala 86:24]
  wire [39:0] vreg_mdu_io_load_kernel; // @[CNN_FU.scala 86:24]
  wire [63:0] vreg_mdu_io_load_vwidth; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_0; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_1; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_2; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_3; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_4; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_5; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_6; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_7; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_8; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_9; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_10; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_11; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_12; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_13; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_14; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_15; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_16; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_17; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_18; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_19; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_20; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_21; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_22; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_23; // @[CNN_FU.scala 86:24]
  wire [15:0] vreg_mdu_io_data_main_24; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_0; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_1; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_2; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_3; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_4; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_5; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_6; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_7; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_8; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_9; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_10; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_11; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_12; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_13; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_14; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_15; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_16; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_17; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_18; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_19; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_20; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_21; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_22; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_23; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_data_kernel_24; // @[CNN_FU.scala 86:24]
  wire [3:0] vreg_mdu_io_data_kernel_vwidth; // @[CNN_FU.scala 86:24]
  wire [7:0] vreg_mdu_io_select_vwidth; // @[CNN_FU.scala 86:24]
  wire [3:0] vreg_mdu_io_act_vwidth; // @[CNN_FU.scala 86:24]
  wire  conv_mdu_clock; // @[CNN_FU.scala 254:24]
  wire  conv_mdu_reset; // @[CNN_FU.scala 254:24]
  wire  conv_mdu_io_conv_valid; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_0; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_1; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_2; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_3; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_4; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_5; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_6; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_7; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_8; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_9; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_10; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_11; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_12; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_13; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_14; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_15; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_16; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_17; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_18; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_19; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_20; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_21; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_22; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_23; // @[CNN_FU.scala 254:24]
  wire [15:0] conv_mdu_io_data_main_24; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_0; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_1; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_2; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_3; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_4; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_5; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_6; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_7; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_8; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_9; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_10; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_11; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_12; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_13; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_14; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_15; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_16; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_17; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_18; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_19; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_20; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_21; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_22; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_23; // @[CNN_FU.scala 254:24]
  wire [7:0] conv_mdu_io_data_kernel_24; // @[CNN_FU.scala 254:24]
  wire [3:0] conv_mdu_io_data_kernel_vwidth; // @[CNN_FU.scala 254:24]
  wire [63:0] conv_mdu_io_conv_res; // @[CNN_FU.scala 254:24]
  wire  conv_mdu_io_conv_ok; // @[CNN_FU.scala 254:24]
  wire [3:0] pool_mdu_io_k; // @[CNN_FU.scala 265:24]
  wire [1:0] pool_mdu_io_agm; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_0; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_1; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_2; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_3; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_4; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_5; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_6; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_7; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_8; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_9; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_10; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_11; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_12; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_13; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_14; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_15; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_16; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_17; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_18; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_19; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_20; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_21; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_22; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_23; // @[CNN_FU.scala 265:24]
  wire [15:0] pool_mdu_io_data_main_24; // @[CNN_FU.scala 265:24]
  wire [63:0] pool_mdu_io_pool_res; // @[CNN_FU.scala 265:24]
  wire [63:0] act_mdu_io_data_main; // @[CNN_FU.scala 275:23]
  wire [63:0] act_mdu_io_data_zero; // @[CNN_FU.scala 275:23]
  wire [3:0] act_mdu_io_data_vwidth; // @[CNN_FU.scala 275:23]
  wire [63:0] act_mdu_io_act_res; // @[CNN_FU.scala 275:23]
  wire  _T_1 = ~io_in_bits_func[3]; // @[CNN_FU.scala 21:27]
  wire  _T_3 = _T_1 & io_in_bits_func[0]; // @[CNN_FU.scala 22:40]
  wire  isConv = _T_3 & io_in_valid; // @[CNN_FU.scala 78:41]
  wire  _T_7 = _T_1 & io_in_bits_func[1]; // @[CNN_FU.scala 23:40]
  wire  isPool = _T_7 & io_in_valid; // @[CNN_FU.scala 79:41]
  wire  _T_11 = _T_1 & io_in_bits_func[2]; // @[CNN_FU.scala 24:40]
  wire  isAct = _T_11 & io_in_valid; // @[CNN_FU.scala 80:41]
  wire  _T_14 = io_in_bits_func[3] & io_in_bits_func[2]; // @[CNN_FU.scala 25:43]
  wire  isLoadD = _T_14 & io_in_valid; // @[CNN_FU.scala 81:41]
  wire  _T_17 = io_in_bits_func[3] & io_in_bits_func[1]; // @[CNN_FU.scala 26:43]
  wire  isLoadP = _T_17 & io_in_valid; // @[CNN_FU.scala 82:41]
  wire  _T_20 = io_in_bits_func[3] & io_in_bits_func[0]; // @[CNN_FU.scala 27:43]
  wire  isLoadW = _T_20 & io_in_valid; // @[CNN_FU.scala 83:41]
  wire  vtype = io_vec_addr[4]; // @[CNN_FU.scala 89:26]
  wire  _T_22 = ~vtype; // @[CNN_FU.scala 90:44]
  wire  isInt16 = vreg_mdu_io_select_vwidth[7] & ~vtype; // @[CNN_FU.scala 90:34]
  wire  isInt8 = vreg_mdu_io_select_vwidth[6] & _T_22 | vreg_mdu_io_select_vwidth[3] & vtype; // @[CNN_FU.scala 91:52]
  wire  isInt4 = vreg_mdu_io_select_vwidth[5] & _T_22 | vreg_mdu_io_select_vwidth[2] & vtype; // @[CNN_FU.scala 92:52]
  wire  isInt2 = vreg_mdu_io_select_vwidth[4] & _T_22 | vreg_mdu_io_select_vwidth[1] & vtype; // @[CNN_FU.scala 93:52]
  wire  isInt1 = vreg_mdu_io_select_vwidth[0] & vtype; // @[CNN_FU.scala 94:33]
  wire [1:0] _T_49 = vreg_mdu_io_select_vwidth[4] + vreg_mdu_io_select_vwidth[5]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_51 = vreg_mdu_io_select_vwidth[6] + vreg_mdu_io_select_vwidth[7]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_53 = _T_49 + _T_51; // @[Bitwise.scala 47:55]
  wire [1:0] _T_63 = vreg_mdu_io_select_vwidth[0] + vreg_mdu_io_select_vwidth[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_65 = vreg_mdu_io_select_vwidth[2] + vreg_mdu_io_select_vwidth[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_67 = _T_63 + _T_65; // @[Bitwise.scala 47:55]
  wire  vwidth_valid = _T_22 & _T_53 == 3'h1 | vtype & _T_67 == 3'h1; // @[CNN_FU.scala 95:80]
  wire  k_valid = io_length_k != 4'h0; // @[CNN_FU.scala 96:30]
  wire [4:0] intNumVec = {isInt16,isInt8,isInt4,isInt2,isInt1}; // @[Cat.scala 30:58]
  reg  state; // @[CNN_FU.scala 105:22]
  reg [63:0] data_stage1_reg; // @[CNN_FU.scala 106:32]
  wire [63:0] int16_src1 = {io_in_bits_src1[63:3],3'h0}; // @[Cat.scala 30:58]
  wire [63:0] int16_src2 = state ? 64'h8 : 64'h0; // @[CNN_FU.scala 112:23]
  wire [2:0] _GEN_5 = {{1'd0}, io_in_bits_src1[2:1]}; // @[CNN_FU.scala 114:39]
  wire [3:0] _T_84 = _GEN_5 + io_length_k[2:0]; // @[CNN_FU.scala 114:39]
  wire  int16_stage2_valid = _T_84 >= 4'h5; // @[CNN_FU.scala 114:60]
  wire [63:0] int8_src2_stage1 = io_in_bits_src1[2] ? 64'h4 : 64'h0; // @[CNN_FU.scala 117:29]
  wire [63:0] int8_src2 = state ? 64'h8 : int8_src2_stage1; // @[CNN_FU.scala 119:22]
  wire [2:0] _T_92 = io_in_bits_src1[2] ? 3'h6 : 3'h3; // @[CNN_FU.scala 120:61]
  wire [2:0] int8_func = state ? 3'h6 : _T_92; // @[CNN_FU.scala 120:22]
  wire [3:0] _T_95 = io_in_bits_src1[2:0] + io_length_k[2:0]; // @[CNN_FU.scala 121:38]
  wire  int8_stage2_valid = _T_95 >= 4'h9; // @[CNN_FU.scala 121:59]
  wire [63:0] int4_src1 = {1'h0,io_in_bits_src1[63:3],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] int4_src2_stage1 = io_in_bits_src1[2] ? 64'h2 : 64'h0; // @[CNN_FU.scala 124:29]
  wire [63:0] int4_src2 = state ? 64'h4 : int4_src2_stage1; // @[CNN_FU.scala 126:22]
  wire [2:0] _T_104 = io_in_bits_src1[2] ? 3'h5 : 3'h6; // @[CNN_FU.scala 127:61]
  wire [2:0] int4_func = state ? 3'h5 : _T_104; // @[CNN_FU.scala 127:22]
  wire [63:0] int2_src1 = {2'h0,io_in_bits_src1[63:3],1'h0}; // @[Cat.scala 30:58]
  wire [63:0] int2_src2_stage1 = io_in_bits_src1[2] ? 64'h1 : 64'h0; // @[CNN_FU.scala 131:29]
  wire [63:0] int2_src2 = state ? 64'h2 : int2_src2_stage1; // @[CNN_FU.scala 133:22]
  wire [2:0] _T_116 = io_in_bits_src1[2] ? 3'h4 : 3'h5; // @[CNN_FU.scala 134:61]
  wire [2:0] int2_func = state ? 3'h4 : _T_116; // @[CNN_FU.scala 134:22]
  wire [63:0] int1_src1 = {3'h0,io_in_bits_src1[63:3]}; // @[Cat.scala 30:58]
  wire [63:0] int1_src2 = state ? 64'h1 : 64'h0; // @[CNN_FU.scala 140:22]
  wire [63:0] _T_126 = 5'h10 == intNumVec ? int16_src1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_128 = 5'h8 == intNumVec ? int16_src1 : _T_126; // @[Mux.scala 80:57]
  wire [63:0] _T_130 = 5'h4 == intNumVec ? int4_src1 : _T_128; // @[Mux.scala 80:57]
  wire [63:0] _T_132 = 5'h2 == intNumVec ? int2_src1 : _T_130; // @[Mux.scala 80:57]
  wire [63:0] loadv_src1 = 5'h1 == intNumVec ? int1_src1 : _T_132; // @[Mux.scala 80:57]
  wire [63:0] _T_135 = 5'h10 == intNumVec ? int16_src2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_137 = 5'h8 == intNumVec ? int8_src2 : _T_135; // @[Mux.scala 80:57]
  wire [63:0] _T_139 = 5'h4 == intNumVec ? int4_src2 : _T_137; // @[Mux.scala 80:57]
  wire [63:0] _T_141 = 5'h2 == intNumVec ? int2_src2 : _T_139; // @[Mux.scala 80:57]
  wire [63:0] loadv_src2 = 5'h1 == intNumVec ? int1_src2 : _T_141; // @[Mux.scala 80:57]
  wire [6:0] _T_144 = 5'h10 == intNumVec ? 7'h3 : 7'h0; // @[Mux.scala 80:57]
  wire [6:0] _T_146 = 5'h8 == intNumVec ? {{4'd0}, int8_func} : _T_144; // @[Mux.scala 80:57]
  wire [6:0] _T_148 = 5'h4 == intNumVec ? {{4'd0}, int4_func} : _T_146; // @[Mux.scala 80:57]
  wire [6:0] _T_150 = 5'h2 == intNumVec ? {{4'd0}, int2_func} : _T_148; // @[Mux.scala 80:57]
  wire [6:0] loadv_func = 5'h1 == intNumVec ? 7'h4 : _T_150; // @[Mux.scala 80:57]
  wire  _T_155 = 5'h8 == intNumVec ? int8_stage2_valid : 5'h10 == intNumVec & int16_stage2_valid; // @[Mux.scala 80:57]
  wire  _T_157 = 5'h4 == intNumVec ? int8_stage2_valid : _T_155; // @[Mux.scala 80:57]
  wire  _T_159 = 5'h2 == intNumVec ? int8_stage2_valid : _T_157; // @[Mux.scala 80:57]
  wire  stage2_valid = 5'h1 == intNumVec ? int8_stage2_valid : _T_159; // @[Mux.scala 80:57]
  wire  _T_161 = ~state; // @[CNN_FU.scala 158:18]
  wire  _T_162 = isLoadD | isLoadP; // @[CNN_FU.scala 160:23]
  wire  _T_165 = ~io_loadv_load_exception; // @[CNN_FU.scala 160:67]
  wire  _GEN_0 = (isLoadD | isLoadP) & stage2_valid & io_loadv_load_valid & ~io_loadv_load_exception | state; // @[CNN_FU.scala 105:22 160:{77,85}]
  wire [63:0] data_stage1 = stage2_valid ? data_stage1_reg : io_loadv_load_data; // @[CNN_FU.scala 169:24]
  wire [79:0] _T_177 = {io_loadv_load_data[15:0],data_stage1}; // @[Cat.scala 30:58]
  wire [79:0] _T_180 = {io_loadv_load_data[31:0],data_stage1[63:16]}; // @[Cat.scala 30:58]
  wire [79:0] _T_183 = {io_loadv_load_data[47:0],data_stage1[63:32]}; // @[Cat.scala 30:58]
  wire [79:0] _T_185 = {io_loadv_load_data,data_stage1[63:48]}; // @[Cat.scala 30:58]
  wire  _T_186 = 2'h0 == io_in_bits_src1[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_187 = 2'h1 == io_in_bits_src1[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_188 = 2'h2 == io_in_bits_src1[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_189 = 2'h3 == io_in_bits_src1[2:1]; // @[LookupTree.scala 24:34]
  wire [79:0] _T_190 = _T_186 ? _T_177 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_191 = _T_187 ? _T_180 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_192 = _T_188 ? _T_183 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_193 = _T_189 ? _T_185 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_194 = _T_190 | _T_191; // @[Mux.scala 27:72]
  wire [79:0] _T_195 = _T_194 | _T_192; // @[Mux.scala 27:72]
  wire [79:0] int16_load_data = _T_195 | _T_193; // @[Mux.scala 27:72]
  wire [7:0] _T_201 = io_loadv_load_data[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_202 = {_T_201,io_loadv_load_data[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_203 = {8'h0,io_loadv_load_data[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_204 = vtype ? _T_202 : _T_203; // @[CNN_FU.scala 38:8]
  wire [7:0] _T_208 = io_loadv_load_data[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_209 = {_T_208,io_loadv_load_data[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_210 = {8'h0,io_loadv_load_data[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_211 = vtype ? _T_209 : _T_210; // @[CNN_FU.scala 38:8]
  wire [7:0] _T_215 = io_loadv_load_data[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_216 = {_T_215,io_loadv_load_data[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_217 = {8'h0,io_loadv_load_data[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_218 = vtype ? _T_216 : _T_217; // @[CNN_FU.scala 38:8]
  wire [7:0] _T_222 = io_loadv_load_data[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_223 = {_T_222,io_loadv_load_data[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_224 = {8'h0,io_loadv_load_data[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_225 = vtype ? _T_223 : _T_224; // @[CNN_FU.scala 38:8]
  wire [7:0] _T_229 = io_loadv_load_data[39] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_230 = {_T_229,io_loadv_load_data[39:32]}; // @[Cat.scala 30:58]
  wire [15:0] _T_231 = {8'h0,io_loadv_load_data[39:32]}; // @[Cat.scala 30:58]
  wire [15:0] _T_232 = vtype ? _T_230 : _T_231; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_233 = {_T_232,_T_225,_T_218,_T_211,_T_204}; // @[Cat.scala 30:58]
  wire [7:0] _T_265 = io_loadv_load_data[47] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_266 = {_T_265,io_loadv_load_data[47:40]}; // @[Cat.scala 30:58]
  wire [15:0] _T_267 = {8'h0,io_loadv_load_data[47:40]}; // @[Cat.scala 30:58]
  wire [15:0] _T_268 = vtype ? _T_266 : _T_267; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_269 = {_T_268,_T_232,_T_225,_T_218,_T_211}; // @[Cat.scala 30:58]
  wire [7:0] _T_301 = io_loadv_load_data[55] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_302 = {_T_301,io_loadv_load_data[55:48]}; // @[Cat.scala 30:58]
  wire [15:0] _T_303 = {8'h0,io_loadv_load_data[55:48]}; // @[Cat.scala 30:58]
  wire [15:0] _T_304 = vtype ? _T_302 : _T_303; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_305 = {_T_304,_T_268,_T_232,_T_225,_T_218}; // @[Cat.scala 30:58]
  wire [7:0] _T_337 = io_loadv_load_data[63] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_338 = {_T_337,io_loadv_load_data[63:56]}; // @[Cat.scala 30:58]
  wire [15:0] _T_339 = {8'h0,io_loadv_load_data[63:56]}; // @[Cat.scala 30:58]
  wire [15:0] _T_340 = vtype ? _T_338 : _T_339; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_341 = {_T_340,_T_304,_T_268,_T_232,_T_225}; // @[Cat.scala 30:58]
  wire [7:0] _T_345 = data_stage1[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_346 = {_T_345,data_stage1[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_347 = {8'h0,data_stage1[7:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_348 = vtype ? _T_346 : _T_347; // @[CNN_FU.scala 38:8]
  wire [7:0] _T_352 = data_stage1[15] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_353 = {_T_352,data_stage1[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_354 = {8'h0,data_stage1[15:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_355 = vtype ? _T_353 : _T_354; // @[CNN_FU.scala 38:8]
  wire [7:0] _T_359 = data_stage1[23] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_360 = {_T_359,data_stage1[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_361 = {8'h0,data_stage1[23:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_362 = vtype ? _T_360 : _T_361; // @[CNN_FU.scala 38:8]
  wire [7:0] _T_366 = data_stage1[31] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_367 = {_T_366,data_stage1[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_368 = {8'h0,data_stage1[31:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_369 = vtype ? _T_367 : _T_368; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_377 = {_T_204,_T_369,_T_362,_T_355,_T_348}; // @[Cat.scala 30:58]
  wire [79:0] _T_413 = {_T_211,_T_204,_T_369,_T_362,_T_355}; // @[Cat.scala 30:58]
  wire [79:0] _T_449 = {_T_218,_T_211,_T_204,_T_369,_T_362}; // @[Cat.scala 30:58]
  wire [79:0] _T_485 = {_T_225,_T_218,_T_211,_T_204,_T_369}; // @[Cat.scala 30:58]
  wire  _T_486 = 3'h0 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_487 = 3'h1 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_488 = 3'h2 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_489 = 3'h3 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_490 = 3'h4 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_491 = 3'h5 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_492 = 3'h6 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_493 = 3'h7 == io_in_bits_src1[2:0]; // @[LookupTree.scala 24:34]
  wire [79:0] _T_494 = _T_486 ? _T_233 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_495 = _T_487 ? _T_269 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_496 = _T_488 ? _T_305 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_497 = _T_489 ? _T_341 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_498 = _T_490 ? _T_377 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_499 = _T_491 ? _T_413 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_500 = _T_492 ? _T_449 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_501 = _T_493 ? _T_485 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_502 = _T_494 | _T_495; // @[Mux.scala 27:72]
  wire [79:0] _T_503 = _T_502 | _T_496; // @[Mux.scala 27:72]
  wire [79:0] _T_504 = _T_503 | _T_497; // @[Mux.scala 27:72]
  wire [79:0] _T_505 = _T_504 | _T_498; // @[Mux.scala 27:72]
  wire [79:0] _T_506 = _T_505 | _T_499; // @[Mux.scala 27:72]
  wire [79:0] _T_507 = _T_506 | _T_500; // @[Mux.scala 27:72]
  wire [79:0] int8_load_data = _T_507 | _T_501; // @[Mux.scala 27:72]
  wire [11:0] _T_513 = io_loadv_load_data[3] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_514 = {_T_513,io_loadv_load_data[3:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_515 = {12'h0,io_loadv_load_data[3:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_516 = vtype ? _T_514 : _T_515; // @[CNN_FU.scala 38:8]
  wire [11:0] _T_520 = io_loadv_load_data[7] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_521 = {_T_520,io_loadv_load_data[7:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_522 = {12'h0,io_loadv_load_data[7:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_523 = vtype ? _T_521 : _T_522; // @[CNN_FU.scala 38:8]
  wire [11:0] _T_527 = io_loadv_load_data[11] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_528 = {_T_527,io_loadv_load_data[11:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_529 = {12'h0,io_loadv_load_data[11:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_530 = vtype ? _T_528 : _T_529; // @[CNN_FU.scala 38:8]
  wire [11:0] _T_534 = io_loadv_load_data[15] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_535 = {_T_534,io_loadv_load_data[15:12]}; // @[Cat.scala 30:58]
  wire [15:0] _T_536 = {12'h0,io_loadv_load_data[15:12]}; // @[Cat.scala 30:58]
  wire [15:0] _T_537 = vtype ? _T_535 : _T_536; // @[CNN_FU.scala 38:8]
  wire [11:0] _T_541 = io_loadv_load_data[19] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_542 = {_T_541,io_loadv_load_data[19:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_543 = {12'h0,io_loadv_load_data[19:16]}; // @[Cat.scala 30:58]
  wire [15:0] _T_544 = vtype ? _T_542 : _T_543; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_545 = {_T_544,_T_537,_T_530,_T_523,_T_516}; // @[Cat.scala 30:58]
  wire [11:0] _T_577 = io_loadv_load_data[23] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_578 = {_T_577,io_loadv_load_data[23:20]}; // @[Cat.scala 30:58]
  wire [15:0] _T_579 = {12'h0,io_loadv_load_data[23:20]}; // @[Cat.scala 30:58]
  wire [15:0] _T_580 = vtype ? _T_578 : _T_579; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_581 = {_T_580,_T_544,_T_537,_T_530,_T_523}; // @[Cat.scala 30:58]
  wire [11:0] _T_613 = io_loadv_load_data[27] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_614 = {_T_613,io_loadv_load_data[27:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_615 = {12'h0,io_loadv_load_data[27:24]}; // @[Cat.scala 30:58]
  wire [15:0] _T_616 = vtype ? _T_614 : _T_615; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_617 = {_T_616,_T_580,_T_544,_T_537,_T_530}; // @[Cat.scala 30:58]
  wire [11:0] _T_649 = io_loadv_load_data[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_650 = {_T_649,io_loadv_load_data[31:28]}; // @[Cat.scala 30:58]
  wire [15:0] _T_651 = {12'h0,io_loadv_load_data[31:28]}; // @[Cat.scala 30:58]
  wire [15:0] _T_652 = vtype ? _T_650 : _T_651; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_653 = {_T_652,_T_616,_T_580,_T_544,_T_537}; // @[Cat.scala 30:58]
  wire [11:0] _T_657 = data_stage1[3] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_658 = {_T_657,data_stage1[3:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_659 = {12'h0,data_stage1[3:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_660 = vtype ? _T_658 : _T_659; // @[CNN_FU.scala 38:8]
  wire [11:0] _T_664 = data_stage1[7] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_665 = {_T_664,data_stage1[7:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_666 = {12'h0,data_stage1[7:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_667 = vtype ? _T_665 : _T_666; // @[CNN_FU.scala 38:8]
  wire [11:0] _T_671 = data_stage1[11] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_672 = {_T_671,data_stage1[11:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_673 = {12'h0,data_stage1[11:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_674 = vtype ? _T_672 : _T_673; // @[CNN_FU.scala 38:8]
  wire [11:0] _T_678 = data_stage1[15] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_679 = {_T_678,data_stage1[15:12]}; // @[Cat.scala 30:58]
  wire [15:0] _T_680 = {12'h0,data_stage1[15:12]}; // @[Cat.scala 30:58]
  wire [15:0] _T_681 = vtype ? _T_679 : _T_680; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_689 = {_T_516,_T_681,_T_674,_T_667,_T_660}; // @[Cat.scala 30:58]
  wire [79:0] _T_725 = {_T_523,_T_516,_T_681,_T_674,_T_667}; // @[Cat.scala 30:58]
  wire [79:0] _T_761 = {_T_530,_T_523,_T_516,_T_681,_T_674}; // @[Cat.scala 30:58]
  wire [79:0] _T_797 = {_T_537,_T_530,_T_523,_T_516,_T_681}; // @[Cat.scala 30:58]
  wire [79:0] _T_806 = _T_486 ? _T_545 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_807 = _T_487 ? _T_581 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_808 = _T_488 ? _T_617 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_809 = _T_489 ? _T_653 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_810 = _T_490 ? _T_689 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_811 = _T_491 ? _T_725 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_812 = _T_492 ? _T_761 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_813 = _T_493 ? _T_797 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_814 = _T_806 | _T_807; // @[Mux.scala 27:72]
  wire [79:0] _T_815 = _T_814 | _T_808; // @[Mux.scala 27:72]
  wire [79:0] _T_816 = _T_815 | _T_809; // @[Mux.scala 27:72]
  wire [79:0] _T_817 = _T_816 | _T_810; // @[Mux.scala 27:72]
  wire [79:0] _T_818 = _T_817 | _T_811; // @[Mux.scala 27:72]
  wire [79:0] _T_819 = _T_818 | _T_812; // @[Mux.scala 27:72]
  wire [79:0] int4_load_data = _T_819 | _T_813; // @[Mux.scala 27:72]
  wire [13:0] _T_825 = io_loadv_load_data[1] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_826 = {_T_825,io_loadv_load_data[1:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_827 = {14'h0,io_loadv_load_data[1:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_828 = vtype ? _T_826 : _T_827; // @[CNN_FU.scala 38:8]
  wire [13:0] _T_832 = io_loadv_load_data[3] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_833 = {_T_832,io_loadv_load_data[3:2]}; // @[Cat.scala 30:58]
  wire [15:0] _T_834 = {14'h0,io_loadv_load_data[3:2]}; // @[Cat.scala 30:58]
  wire [15:0] _T_835 = vtype ? _T_833 : _T_834; // @[CNN_FU.scala 38:8]
  wire [13:0] _T_839 = io_loadv_load_data[5] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_840 = {_T_839,io_loadv_load_data[5:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_841 = {14'h0,io_loadv_load_data[5:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_842 = vtype ? _T_840 : _T_841; // @[CNN_FU.scala 38:8]
  wire [13:0] _T_846 = io_loadv_load_data[7] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_847 = {_T_846,io_loadv_load_data[7:6]}; // @[Cat.scala 30:58]
  wire [15:0] _T_848 = {14'h0,io_loadv_load_data[7:6]}; // @[Cat.scala 30:58]
  wire [15:0] _T_849 = vtype ? _T_847 : _T_848; // @[CNN_FU.scala 38:8]
  wire [13:0] _T_853 = io_loadv_load_data[9] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_854 = {_T_853,io_loadv_load_data[9:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_855 = {14'h0,io_loadv_load_data[9:8]}; // @[Cat.scala 30:58]
  wire [15:0] _T_856 = vtype ? _T_854 : _T_855; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_857 = {_T_856,_T_849,_T_842,_T_835,_T_828}; // @[Cat.scala 30:58]
  wire [13:0] _T_889 = io_loadv_load_data[11] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_890 = {_T_889,io_loadv_load_data[11:10]}; // @[Cat.scala 30:58]
  wire [15:0] _T_891 = {14'h0,io_loadv_load_data[11:10]}; // @[Cat.scala 30:58]
  wire [15:0] _T_892 = vtype ? _T_890 : _T_891; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_893 = {_T_892,_T_856,_T_849,_T_842,_T_835}; // @[Cat.scala 30:58]
  wire [13:0] _T_925 = io_loadv_load_data[13] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_926 = {_T_925,io_loadv_load_data[13:12]}; // @[Cat.scala 30:58]
  wire [15:0] _T_927 = {14'h0,io_loadv_load_data[13:12]}; // @[Cat.scala 30:58]
  wire [15:0] _T_928 = vtype ? _T_926 : _T_927; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_929 = {_T_928,_T_892,_T_856,_T_849,_T_842}; // @[Cat.scala 30:58]
  wire [13:0] _T_961 = io_loadv_load_data[15] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_962 = {_T_961,io_loadv_load_data[15:14]}; // @[Cat.scala 30:58]
  wire [15:0] _T_963 = {14'h0,io_loadv_load_data[15:14]}; // @[Cat.scala 30:58]
  wire [15:0] _T_964 = vtype ? _T_962 : _T_963; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_965 = {_T_964,_T_928,_T_892,_T_856,_T_849}; // @[Cat.scala 30:58]
  wire [13:0] _T_969 = data_stage1[1] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_970 = {_T_969,data_stage1[1:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_971 = {14'h0,data_stage1[1:0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_972 = vtype ? _T_970 : _T_971; // @[CNN_FU.scala 38:8]
  wire [13:0] _T_976 = data_stage1[3] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_977 = {_T_976,data_stage1[3:2]}; // @[Cat.scala 30:58]
  wire [15:0] _T_978 = {14'h0,data_stage1[3:2]}; // @[Cat.scala 30:58]
  wire [15:0] _T_979 = vtype ? _T_977 : _T_978; // @[CNN_FU.scala 38:8]
  wire [13:0] _T_983 = data_stage1[5] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_984 = {_T_983,data_stage1[5:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_985 = {14'h0,data_stage1[5:4]}; // @[Cat.scala 30:58]
  wire [15:0] _T_986 = vtype ? _T_984 : _T_985; // @[CNN_FU.scala 38:8]
  wire [13:0] _T_990 = data_stage1[7] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_991 = {_T_990,data_stage1[7:6]}; // @[Cat.scala 30:58]
  wire [15:0] _T_992 = {14'h0,data_stage1[7:6]}; // @[Cat.scala 30:58]
  wire [15:0] _T_993 = vtype ? _T_991 : _T_992; // @[CNN_FU.scala 38:8]
  wire [79:0] _T_1001 = {_T_828,_T_993,_T_986,_T_979,_T_972}; // @[Cat.scala 30:58]
  wire [79:0] _T_1037 = {_T_835,_T_828,_T_993,_T_986,_T_979}; // @[Cat.scala 30:58]
  wire [79:0] _T_1073 = {_T_842,_T_835,_T_828,_T_993,_T_986}; // @[Cat.scala 30:58]
  wire [79:0] _T_1109 = {_T_849,_T_842,_T_835,_T_828,_T_993}; // @[Cat.scala 30:58]
  wire [79:0] _T_1118 = _T_486 ? _T_857 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1119 = _T_487 ? _T_893 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1120 = _T_488 ? _T_929 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1121 = _T_489 ? _T_965 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1122 = _T_490 ? _T_1001 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1123 = _T_491 ? _T_1037 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1124 = _T_492 ? _T_1073 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1125 = _T_493 ? _T_1109 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1126 = _T_1118 | _T_1119; // @[Mux.scala 27:72]
  wire [79:0] _T_1127 = _T_1126 | _T_1120; // @[Mux.scala 27:72]
  wire [79:0] _T_1128 = _T_1127 | _T_1121; // @[Mux.scala 27:72]
  wire [79:0] _T_1129 = _T_1128 | _T_1122; // @[Mux.scala 27:72]
  wire [79:0] _T_1130 = _T_1129 | _T_1123; // @[Mux.scala 27:72]
  wire [79:0] _T_1131 = _T_1130 | _T_1124; // @[Mux.scala 27:72]
  wire [79:0] int2_load_data = _T_1131 | _T_1125; // @[Mux.scala 27:72]
  wire [79:0] _T_1144 = {15'h0,io_loadv_load_data[4],15'h0,io_loadv_load_data[3],15'h0,io_loadv_load_data[2],15'h0,
    io_loadv_load_data[1],15'h0,io_loadv_load_data[0]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1155 = {15'h0,io_loadv_load_data[5],15'h0,io_loadv_load_data[4],15'h0,io_loadv_load_data[3],15'h0,
    io_loadv_load_data[2],15'h0,io_loadv_load_data[1]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1166 = {15'h0,io_loadv_load_data[6],15'h0,io_loadv_load_data[5],15'h0,io_loadv_load_data[4],15'h0,
    io_loadv_load_data[3],15'h0,io_loadv_load_data[2]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1177 = {15'h0,io_loadv_load_data[7],15'h0,io_loadv_load_data[6],15'h0,io_loadv_load_data[5],15'h0,
    io_loadv_load_data[4],15'h0,io_loadv_load_data[3]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1188 = {15'h0,io_loadv_load_data[0],15'h0,data_stage1[7],15'h0,data_stage1[6],15'h0,data_stage1[5],15'h0
    ,data_stage1[4]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1199 = {15'h0,io_loadv_load_data[1],15'h0,io_loadv_load_data[0],15'h0,data_stage1[7],15'h0,data_stage1[
    6],15'h0,data_stage1[5]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1210 = {15'h0,io_loadv_load_data[2],15'h0,io_loadv_load_data[1],15'h0,io_loadv_load_data[0],15'h0,
    data_stage1[7],15'h0,data_stage1[6]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1221 = {15'h0,io_loadv_load_data[3],15'h0,io_loadv_load_data[2],15'h0,io_loadv_load_data[1],15'h0,
    io_loadv_load_data[0],15'h0,data_stage1[7]}; // @[Cat.scala 30:58]
  wire [79:0] _T_1230 = _T_486 ? _T_1144 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1231 = _T_487 ? _T_1155 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1232 = _T_488 ? _T_1166 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1233 = _T_489 ? _T_1177 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1234 = _T_490 ? _T_1188 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1235 = _T_491 ? _T_1199 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1236 = _T_492 ? _T_1210 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1237 = _T_493 ? _T_1221 : 80'h0; // @[Mux.scala 27:72]
  wire [79:0] _T_1238 = _T_1230 | _T_1231; // @[Mux.scala 27:72]
  wire [79:0] _T_1239 = _T_1238 | _T_1232; // @[Mux.scala 27:72]
  wire [79:0] _T_1240 = _T_1239 | _T_1233; // @[Mux.scala 27:72]
  wire [79:0] _T_1241 = _T_1240 | _T_1234; // @[Mux.scala 27:72]
  wire [79:0] _T_1242 = _T_1241 | _T_1235; // @[Mux.scala 27:72]
  wire [79:0] _T_1243 = _T_1242 | _T_1236; // @[Mux.scala 27:72]
  wire [79:0] int1_load_data = _T_1243 | _T_1237; // @[Mux.scala 27:72]
  wire [79:0] _T_1246 = 5'h10 == intNumVec ? int16_load_data : 80'h0; // @[Mux.scala 80:57]
  wire [79:0] _T_1248 = 5'h8 == intNumVec ? int8_load_data : _T_1246; // @[Mux.scala 80:57]
  wire [79:0] _T_1250 = 5'h4 == intNumVec ? int4_load_data : _T_1248; // @[Mux.scala 80:57]
  wire [79:0] _T_1252 = 5'h2 == intNumVec ? int2_load_data : _T_1250; // @[Mux.scala 80:57]
  wire [79:0] loadv_data = 5'h1 == intNumVec ? int1_load_data : _T_1252; // @[Mux.scala 80:57]
  wire [15:0] loadv_data_elem_0 = io_length_k[2:0] >= 3'h1 ? loadv_data[15:0] : 16'h0; // @[CNN_FU.scala 229:30]
  wire [15:0] loadv_data_elem_1 = io_length_k[2:0] >= 3'h2 ? loadv_data[31:16] : 16'h0; // @[CNN_FU.scala 229:30]
  wire [15:0] loadv_data_elem_2 = io_length_k[2:0] >= 3'h3 ? loadv_data[47:32] : 16'h0; // @[CNN_FU.scala 229:30]
  wire [15:0] loadv_data_elem_3 = io_length_k[2:0] >= 3'h4 ? loadv_data[63:48] : 16'h0; // @[CNN_FU.scala 229:30]
  wire [15:0] loadv_data_elem_4 = io_length_k[2:0] >= 3'h5 ? loadv_data[79:64] : 16'h0; // @[CNN_FU.scala 229:30]
  wire [63:0] _T_1276 = {loadv_data_elem_3,loadv_data_elem_2,loadv_data_elem_1,loadv_data_elem_0}; // @[Cat.scala 30:58]
  wire [31:0] _T_1284 = {loadv_data_elem_3[7:0],loadv_data_elem_2[7:0],loadv_data_elem_1[7:0],loadv_data_elem_0[7:0]}; // @[Cat.scala 30:58]
  wire  loadv_valid = stage2_valid ? state & io_loadv_load_valid | _T_161 & io_loadv_load_valid &
    io_loadv_load_exception : io_loadv_load_valid; // @[CNN_FU.scala 234:24]
  wire  _T_1293 = _T_162 & vwidth_valid & k_valid; // @[CNN_FU.scala 236:58]
  wire  _T_1294 = _T_162 & vwidth_valid & k_valid | isLoadW; // @[CNN_FU.scala 236:69]
  wire  _T_1304 = _T_1293 ? loadv_valid : 1'h1; // @[CNN_FU.scala 240:45]
  wire  lv_valid = isLoadW ? io_loadv_load_valid : _T_1304; // @[CNN_FU.scala 240:21]
  wire  _T_1313 = isConv ? conv_mdu_io_conv_ok : lv_valid; // @[CNN_FU.scala 284:77]
  wire [63:0] _T_1317 = isPool ? pool_mdu_io_pool_res : conv_mdu_io_conv_res; // @[CNN_FU.scala 285:41]
  CNNVectorRegFile vreg_mdu ( // @[CNN_FU.scala 86:24]
    .clock(vreg_mdu_clock),
    .io_vaddr(vreg_mdu_io_vaddr),
    .io_vtag(vreg_mdu_io_vtag),
    .io_vop(vreg_mdu_io_vop),
    .io_k(vreg_mdu_io_k),
    .io_vwen(vreg_mdu_io_vwen),
    .io_load_data(vreg_mdu_io_load_data),
    .io_load_kernel(vreg_mdu_io_load_kernel),
    .io_load_vwidth(vreg_mdu_io_load_vwidth),
    .io_data_main_0(vreg_mdu_io_data_main_0),
    .io_data_main_1(vreg_mdu_io_data_main_1),
    .io_data_main_2(vreg_mdu_io_data_main_2),
    .io_data_main_3(vreg_mdu_io_data_main_3),
    .io_data_main_4(vreg_mdu_io_data_main_4),
    .io_data_main_5(vreg_mdu_io_data_main_5),
    .io_data_main_6(vreg_mdu_io_data_main_6),
    .io_data_main_7(vreg_mdu_io_data_main_7),
    .io_data_main_8(vreg_mdu_io_data_main_8),
    .io_data_main_9(vreg_mdu_io_data_main_9),
    .io_data_main_10(vreg_mdu_io_data_main_10),
    .io_data_main_11(vreg_mdu_io_data_main_11),
    .io_data_main_12(vreg_mdu_io_data_main_12),
    .io_data_main_13(vreg_mdu_io_data_main_13),
    .io_data_main_14(vreg_mdu_io_data_main_14),
    .io_data_main_15(vreg_mdu_io_data_main_15),
    .io_data_main_16(vreg_mdu_io_data_main_16),
    .io_data_main_17(vreg_mdu_io_data_main_17),
    .io_data_main_18(vreg_mdu_io_data_main_18),
    .io_data_main_19(vreg_mdu_io_data_main_19),
    .io_data_main_20(vreg_mdu_io_data_main_20),
    .io_data_main_21(vreg_mdu_io_data_main_21),
    .io_data_main_22(vreg_mdu_io_data_main_22),
    .io_data_main_23(vreg_mdu_io_data_main_23),
    .io_data_main_24(vreg_mdu_io_data_main_24),
    .io_data_kernel_0(vreg_mdu_io_data_kernel_0),
    .io_data_kernel_1(vreg_mdu_io_data_kernel_1),
    .io_data_kernel_2(vreg_mdu_io_data_kernel_2),
    .io_data_kernel_3(vreg_mdu_io_data_kernel_3),
    .io_data_kernel_4(vreg_mdu_io_data_kernel_4),
    .io_data_kernel_5(vreg_mdu_io_data_kernel_5),
    .io_data_kernel_6(vreg_mdu_io_data_kernel_6),
    .io_data_kernel_7(vreg_mdu_io_data_kernel_7),
    .io_data_kernel_8(vreg_mdu_io_data_kernel_8),
    .io_data_kernel_9(vreg_mdu_io_data_kernel_9),
    .io_data_kernel_10(vreg_mdu_io_data_kernel_10),
    .io_data_kernel_11(vreg_mdu_io_data_kernel_11),
    .io_data_kernel_12(vreg_mdu_io_data_kernel_12),
    .io_data_kernel_13(vreg_mdu_io_data_kernel_13),
    .io_data_kernel_14(vreg_mdu_io_data_kernel_14),
    .io_data_kernel_15(vreg_mdu_io_data_kernel_15),
    .io_data_kernel_16(vreg_mdu_io_data_kernel_16),
    .io_data_kernel_17(vreg_mdu_io_data_kernel_17),
    .io_data_kernel_18(vreg_mdu_io_data_kernel_18),
    .io_data_kernel_19(vreg_mdu_io_data_kernel_19),
    .io_data_kernel_20(vreg_mdu_io_data_kernel_20),
    .io_data_kernel_21(vreg_mdu_io_data_kernel_21),
    .io_data_kernel_22(vreg_mdu_io_data_kernel_22),
    .io_data_kernel_23(vreg_mdu_io_data_kernel_23),
    .io_data_kernel_24(vreg_mdu_io_data_kernel_24),
    .io_data_kernel_vwidth(vreg_mdu_io_data_kernel_vwidth),
    .io_select_vwidth(vreg_mdu_io_select_vwidth),
    .io_act_vwidth(vreg_mdu_io_act_vwidth)
  );
  CNNConv conv_mdu ( // @[CNN_FU.scala 254:24]
    .clock(conv_mdu_clock),
    .reset(conv_mdu_reset),
    .io_conv_valid(conv_mdu_io_conv_valid),
    .io_data_main_0(conv_mdu_io_data_main_0),
    .io_data_main_1(conv_mdu_io_data_main_1),
    .io_data_main_2(conv_mdu_io_data_main_2),
    .io_data_main_3(conv_mdu_io_data_main_3),
    .io_data_main_4(conv_mdu_io_data_main_4),
    .io_data_main_5(conv_mdu_io_data_main_5),
    .io_data_main_6(conv_mdu_io_data_main_6),
    .io_data_main_7(conv_mdu_io_data_main_7),
    .io_data_main_8(conv_mdu_io_data_main_8),
    .io_data_main_9(conv_mdu_io_data_main_9),
    .io_data_main_10(conv_mdu_io_data_main_10),
    .io_data_main_11(conv_mdu_io_data_main_11),
    .io_data_main_12(conv_mdu_io_data_main_12),
    .io_data_main_13(conv_mdu_io_data_main_13),
    .io_data_main_14(conv_mdu_io_data_main_14),
    .io_data_main_15(conv_mdu_io_data_main_15),
    .io_data_main_16(conv_mdu_io_data_main_16),
    .io_data_main_17(conv_mdu_io_data_main_17),
    .io_data_main_18(conv_mdu_io_data_main_18),
    .io_data_main_19(conv_mdu_io_data_main_19),
    .io_data_main_20(conv_mdu_io_data_main_20),
    .io_data_main_21(conv_mdu_io_data_main_21),
    .io_data_main_22(conv_mdu_io_data_main_22),
    .io_data_main_23(conv_mdu_io_data_main_23),
    .io_data_main_24(conv_mdu_io_data_main_24),
    .io_data_kernel_0(conv_mdu_io_data_kernel_0),
    .io_data_kernel_1(conv_mdu_io_data_kernel_1),
    .io_data_kernel_2(conv_mdu_io_data_kernel_2),
    .io_data_kernel_3(conv_mdu_io_data_kernel_3),
    .io_data_kernel_4(conv_mdu_io_data_kernel_4),
    .io_data_kernel_5(conv_mdu_io_data_kernel_5),
    .io_data_kernel_6(conv_mdu_io_data_kernel_6),
    .io_data_kernel_7(conv_mdu_io_data_kernel_7),
    .io_data_kernel_8(conv_mdu_io_data_kernel_8),
    .io_data_kernel_9(conv_mdu_io_data_kernel_9),
    .io_data_kernel_10(conv_mdu_io_data_kernel_10),
    .io_data_kernel_11(conv_mdu_io_data_kernel_11),
    .io_data_kernel_12(conv_mdu_io_data_kernel_12),
    .io_data_kernel_13(conv_mdu_io_data_kernel_13),
    .io_data_kernel_14(conv_mdu_io_data_kernel_14),
    .io_data_kernel_15(conv_mdu_io_data_kernel_15),
    .io_data_kernel_16(conv_mdu_io_data_kernel_16),
    .io_data_kernel_17(conv_mdu_io_data_kernel_17),
    .io_data_kernel_18(conv_mdu_io_data_kernel_18),
    .io_data_kernel_19(conv_mdu_io_data_kernel_19),
    .io_data_kernel_20(conv_mdu_io_data_kernel_20),
    .io_data_kernel_21(conv_mdu_io_data_kernel_21),
    .io_data_kernel_22(conv_mdu_io_data_kernel_22),
    .io_data_kernel_23(conv_mdu_io_data_kernel_23),
    .io_data_kernel_24(conv_mdu_io_data_kernel_24),
    .io_data_kernel_vwidth(conv_mdu_io_data_kernel_vwidth),
    .io_conv_res(conv_mdu_io_conv_res),
    .io_conv_ok(conv_mdu_io_conv_ok)
  );
  CNNPool pool_mdu ( // @[CNN_FU.scala 265:24]
    .io_k(pool_mdu_io_k),
    .io_agm(pool_mdu_io_agm),
    .io_data_main_0(pool_mdu_io_data_main_0),
    .io_data_main_1(pool_mdu_io_data_main_1),
    .io_data_main_2(pool_mdu_io_data_main_2),
    .io_data_main_3(pool_mdu_io_data_main_3),
    .io_data_main_4(pool_mdu_io_data_main_4),
    .io_data_main_5(pool_mdu_io_data_main_5),
    .io_data_main_6(pool_mdu_io_data_main_6),
    .io_data_main_7(pool_mdu_io_data_main_7),
    .io_data_main_8(pool_mdu_io_data_main_8),
    .io_data_main_9(pool_mdu_io_data_main_9),
    .io_data_main_10(pool_mdu_io_data_main_10),
    .io_data_main_11(pool_mdu_io_data_main_11),
    .io_data_main_12(pool_mdu_io_data_main_12),
    .io_data_main_13(pool_mdu_io_data_main_13),
    .io_data_main_14(pool_mdu_io_data_main_14),
    .io_data_main_15(pool_mdu_io_data_main_15),
    .io_data_main_16(pool_mdu_io_data_main_16),
    .io_data_main_17(pool_mdu_io_data_main_17),
    .io_data_main_18(pool_mdu_io_data_main_18),
    .io_data_main_19(pool_mdu_io_data_main_19),
    .io_data_main_20(pool_mdu_io_data_main_20),
    .io_data_main_21(pool_mdu_io_data_main_21),
    .io_data_main_22(pool_mdu_io_data_main_22),
    .io_data_main_23(pool_mdu_io_data_main_23),
    .io_data_main_24(pool_mdu_io_data_main_24),
    .io_pool_res(pool_mdu_io_pool_res)
  );
  CNNAct act_mdu ( // @[CNN_FU.scala 275:23]
    .io_data_main(act_mdu_io_data_main),
    .io_data_zero(act_mdu_io_data_zero),
    .io_data_vwidth(act_mdu_io_data_vwidth),
    .io_act_res(act_mdu_io_act_res)
  );
  assign io_out_valid = io_in_valid & (isAct | (isPool | _T_1313)); // @[CNN_FU.scala 284:25]
  assign io_out_bits = isAct ? act_mdu_io_act_res : _T_1317; // @[CNN_FU.scala 285:21]
  assign io_loadv_valid = _T_162 & vwidth_valid & k_valid | isLoadW; // @[CNN_FU.scala 236:69]
  assign io_loadv_src1 = _T_162 ? loadv_src1 : io_in_bits_src1; // @[CNN_FU.scala 237:23]
  assign io_loadv_src2 = _T_162 ? loadv_src2 : io_imm; // @[CNN_FU.scala 238:23]
  assign io_loadv_func = _T_162 ? loadv_func : 7'h3; // @[CNN_FU.scala 239:23]
  assign vreg_mdu_clock = clock;
  assign vreg_mdu_io_vaddr = io_vec_addr; // @[CNN_FU.scala 244:27]
  assign vreg_mdu_io_vtag = io_vtag; // @[CNN_FU.scala 245:27]
  assign vreg_mdu_io_vop = io_in_bits_func[2:0]; // @[CNN_FU.scala 246:34]
  assign vreg_mdu_io_k = io_length_k; // @[CNN_FU.scala 247:27]
  assign vreg_mdu_io_vwen = lv_valid & _T_1294 & _T_165; // @[CNN_FU.scala 248:103]
  assign vreg_mdu_io_load_data = {loadv_data_elem_4,_T_1276}; // @[Cat.scala 30:58]
  assign vreg_mdu_io_load_kernel = {loadv_data_elem_4[7:0],_T_1284}; // @[Cat.scala 30:58]
  assign vreg_mdu_io_load_vwidth = io_loadv_load_data; // @[CNN_FU.scala 251:27]
  assign conv_mdu_clock = clock;
  assign conv_mdu_reset = reset;
  assign conv_mdu_io_conv_valid = _T_3 & io_in_valid; // @[CNN_FU.scala 78:41]
  assign conv_mdu_io_data_main_0 = vreg_mdu_io_data_main_0; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_1 = vreg_mdu_io_data_main_1; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_2 = vreg_mdu_io_data_main_2; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_3 = vreg_mdu_io_data_main_3; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_4 = vreg_mdu_io_data_main_4; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_5 = vreg_mdu_io_data_main_5; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_6 = vreg_mdu_io_data_main_6; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_7 = vreg_mdu_io_data_main_7; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_8 = vreg_mdu_io_data_main_8; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_9 = vreg_mdu_io_data_main_9; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_10 = vreg_mdu_io_data_main_10; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_11 = vreg_mdu_io_data_main_11; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_12 = vreg_mdu_io_data_main_12; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_13 = vreg_mdu_io_data_main_13; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_14 = vreg_mdu_io_data_main_14; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_15 = vreg_mdu_io_data_main_15; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_16 = vreg_mdu_io_data_main_16; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_17 = vreg_mdu_io_data_main_17; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_18 = vreg_mdu_io_data_main_18; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_19 = vreg_mdu_io_data_main_19; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_20 = vreg_mdu_io_data_main_20; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_21 = vreg_mdu_io_data_main_21; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_22 = vreg_mdu_io_data_main_22; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_23 = vreg_mdu_io_data_main_23; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_main_24 = vreg_mdu_io_data_main_24; // @[CNN_FU.scala 257:34]
  assign conv_mdu_io_data_kernel_0 = vreg_mdu_io_data_kernel_0; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_1 = vreg_mdu_io_data_kernel_1; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_2 = vreg_mdu_io_data_kernel_2; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_3 = vreg_mdu_io_data_kernel_3; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_4 = vreg_mdu_io_data_kernel_4; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_5 = vreg_mdu_io_data_kernel_5; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_6 = vreg_mdu_io_data_kernel_6; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_7 = vreg_mdu_io_data_kernel_7; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_8 = vreg_mdu_io_data_kernel_8; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_9 = vreg_mdu_io_data_kernel_9; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_10 = vreg_mdu_io_data_kernel_10; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_11 = vreg_mdu_io_data_kernel_11; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_12 = vreg_mdu_io_data_kernel_12; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_13 = vreg_mdu_io_data_kernel_13; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_14 = vreg_mdu_io_data_kernel_14; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_15 = vreg_mdu_io_data_kernel_15; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_16 = vreg_mdu_io_data_kernel_16; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_17 = vreg_mdu_io_data_kernel_17; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_18 = vreg_mdu_io_data_kernel_18; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_19 = vreg_mdu_io_data_kernel_19; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_20 = vreg_mdu_io_data_kernel_20; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_21 = vreg_mdu_io_data_kernel_21; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_22 = vreg_mdu_io_data_kernel_22; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_23 = vreg_mdu_io_data_kernel_23; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_24 = vreg_mdu_io_data_kernel_24; // @[CNN_FU.scala 258:34]
  assign conv_mdu_io_data_kernel_vwidth = vreg_mdu_io_data_kernel_vwidth; // @[CNN_FU.scala 260:34]
  assign pool_mdu_io_k = io_length_k; // @[CNN_FU.scala 267:27]
  assign pool_mdu_io_agm = io_algorithm; // @[CNN_FU.scala 268:27]
  assign pool_mdu_io_data_main_0 = vreg_mdu_io_data_main_0; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_1 = vreg_mdu_io_data_main_1; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_2 = vreg_mdu_io_data_main_2; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_3 = vreg_mdu_io_data_main_3; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_4 = vreg_mdu_io_data_main_4; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_5 = vreg_mdu_io_data_main_5; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_6 = vreg_mdu_io_data_main_6; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_7 = vreg_mdu_io_data_main_7; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_8 = vreg_mdu_io_data_main_8; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_9 = vreg_mdu_io_data_main_9; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_10 = vreg_mdu_io_data_main_10; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_11 = vreg_mdu_io_data_main_11; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_12 = vreg_mdu_io_data_main_12; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_13 = vreg_mdu_io_data_main_13; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_14 = vreg_mdu_io_data_main_14; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_15 = vreg_mdu_io_data_main_15; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_16 = vreg_mdu_io_data_main_16; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_17 = vreg_mdu_io_data_main_17; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_18 = vreg_mdu_io_data_main_18; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_19 = vreg_mdu_io_data_main_19; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_20 = vreg_mdu_io_data_main_20; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_21 = vreg_mdu_io_data_main_21; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_22 = vreg_mdu_io_data_main_22; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_23 = vreg_mdu_io_data_main_23; // @[CNN_FU.scala 269:27]
  assign pool_mdu_io_data_main_24 = vreg_mdu_io_data_main_24; // @[CNN_FU.scala 269:27]
  assign act_mdu_io_data_main = io_in_bits_src1; // @[CNN_FU.scala 277:26]
  assign act_mdu_io_data_zero = io_in_bits_src2; // @[CNN_FU.scala 278:26]
  assign act_mdu_io_data_vwidth = vreg_mdu_io_act_vwidth; // @[CNN_FU.scala 279:26]
  always @(posedge clock) begin
    if (reset) begin // @[CNN_FU.scala 105:22]
      state <= 1'h0; // @[CNN_FU.scala 105:22]
    end else if (~state) begin // @[CNN_FU.scala 158:18]
      state <= _GEN_0;
    end else if (state) begin // @[CNN_FU.scala 158:18]
      if (io_loadv_load_valid) begin // @[CNN_FU.scala 163:26]
        state <= 1'h0; // @[CNN_FU.scala 163:34]
      end
    end
    if (reset) begin // @[CNN_FU.scala 106:32]
      data_stage1_reg <= 64'h0; // @[CNN_FU.scala 106:32]
    end else if (_T_161 & _T_162 & stage2_valid & io_loadv_load_valid & _T_165) begin // @[CNN_FU.scala 166:97]
      data_stage1_reg <= io_loadv_load_data; // @[CNN_FU.scala 166:115]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  data_stage1_reg = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__wdata,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  output        io__dmem_resp_ready,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__isMMIO,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  input         DTLBPF,
  input         DTLBENABLE,
  input         ISAMO2,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addrLatch; // @[UnpipelinedLSU.scala 333:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[UnpipelinedLSU.scala 334:23]
  wire  _T_1 = ~isStore; // @[UnpipelinedLSU.scala 335:21]
  wire  partialLoad = ~isStore & io__in_bits_func != 7'h3; // @[UnpipelinedLSU.scala 335:30]
  reg [1:0] state; // @[UnpipelinedLSU.scala 338:22]
  wire  _T_4 = io__dmem_req_ready & io__dmem_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_2 = DTLBFINISH & DTLBPF ? 2'h0 : state; // @[UnpipelinedLSU.scala 338:22 358:{36,44}]
  wire  _T_14 = io__dmem_resp_ready & io__dmem_resp_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_15 = partialLoad ? 2'h3 : 2'h0; // @[UnpipelinedLSU.scala 361:62]
  wire [1:0] _GEN_4 = _T_14 ? _T_15 : state; // @[UnpipelinedLSU.scala 338:22 361:{48,56}]
  wire [1:0] _GEN_5 = 2'h3 == state ? 2'h0 : state; // @[UnpipelinedLSU.scala 351:18 338:22 362:32]
  wire [1:0] size = io__in_bits_func[1:0]; // @[UnpipelinedLSU.scala 369:18]
  wire [63:0] _T_20 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],
    io__wdata[7:0],io__wdata[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_23 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_25 = {io__wdata[31:0],io__wdata[31:0]}; // @[Cat.scala 30:58]
  wire  _T_26 = 2'h0 == size; // @[LookupTree.scala 24:34]
  wire  _T_27 = 2'h1 == size; // @[LookupTree.scala 24:34]
  wire  _T_28 = 2'h2 == size; // @[LookupTree.scala 24:34]
  wire  _T_29 = 2'h3 == size; // @[LookupTree.scala 24:34]
  wire [63:0] _T_30 = _T_26 ? _T_20 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_31 = _T_27 ? _T_23 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_32 = _T_28 ? _T_25 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_33 = _T_29 ? io__wdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_34 = _T_30 | _T_31; // @[Mux.scala 27:72]
  wire [63:0] _T_35 = _T_34 | _T_32; // @[Mux.scala 27:72]
  wire [1:0] _T_42 = _T_27 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_43 = _T_28 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_44 = _T_29 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_13 = {{1'd0}, _T_26}; // @[Mux.scala 27:72]
  wire [1:0] _T_45 = _GEN_13 | _T_42; // @[Mux.scala 27:72]
  wire [3:0] _GEN_14 = {{2'd0}, _T_45}; // @[Mux.scala 27:72]
  wire [3:0] _T_46 = _GEN_14 | _T_43; // @[Mux.scala 27:72]
  wire [7:0] _GEN_15 = {{4'd0}, _T_46}; // @[Mux.scala 27:72]
  wire [7:0] _T_47 = _GEN_15 | _T_44; // @[Mux.scala 27:72]
  wire [14:0] _GEN_23 = {{7'd0}, _T_47}; // @[UnpipelinedLSU.scala 306:8]
  wire [14:0] reqWmask = _GEN_23 << io__in_bits_src1[2:0]; // @[UnpipelinedLSU.scala 306:8]
  wire  _T_64 = partialLoad ? state == 2'h3 : _T_14 & state == 2'h2; // @[UnpipelinedLSU.scala 382:114]
  reg [63:0] rdataLatch; // @[UnpipelinedLSU.scala 388:27]
  wire  _T_77 = 3'h0 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_78 = 3'h1 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_79 = 3'h2 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_80 = 3'h3 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_81 = 3'h4 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_82 = 3'h5 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_83 = 3'h6 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_84 = 3'h7 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_85 = _T_77 ? rdataLatch : 64'h0; // @[Mux.scala 27:72]
  wire [55:0] _T_86 = _T_78 ? rdataLatch[63:8] : 56'h0; // @[Mux.scala 27:72]
  wire [47:0] _T_87 = _T_79 ? rdataLatch[63:16] : 48'h0; // @[Mux.scala 27:72]
  wire [39:0] _T_88 = _T_80 ? rdataLatch[63:24] : 40'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_89 = _T_81 ? rdataLatch[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_90 = _T_82 ? rdataLatch[63:40] : 24'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_91 = _T_83 ? rdataLatch[63:48] : 16'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_92 = _T_84 ? rdataLatch[63:56] : 8'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_16 = {{8'd0}, _T_86}; // @[Mux.scala 27:72]
  wire [63:0] _T_93 = _T_85 | _GEN_16; // @[Mux.scala 27:72]
  wire [63:0] _GEN_17 = {{16'd0}, _T_87}; // @[Mux.scala 27:72]
  wire [63:0] _T_94 = _T_93 | _GEN_17; // @[Mux.scala 27:72]
  wire [63:0] _GEN_18 = {{24'd0}, _T_88}; // @[Mux.scala 27:72]
  wire [63:0] _T_95 = _T_94 | _GEN_18; // @[Mux.scala 27:72]
  wire [63:0] _GEN_19 = {{32'd0}, _T_89}; // @[Mux.scala 27:72]
  wire [63:0] _T_96 = _T_95 | _GEN_19; // @[Mux.scala 27:72]
  wire [63:0] _GEN_20 = {{40'd0}, _T_90}; // @[Mux.scala 27:72]
  wire [63:0] _T_97 = _T_96 | _GEN_20; // @[Mux.scala 27:72]
  wire [63:0] _GEN_21 = {{48'd0}, _T_91}; // @[Mux.scala 27:72]
  wire [63:0] _T_98 = _T_97 | _GEN_21; // @[Mux.scala 27:72]
  wire [63:0] _GEN_22 = {{56'd0}, _T_92}; // @[Mux.scala 27:72]
  wire [63:0] rdataSel = _T_98 | _GEN_22; // @[Mux.scala 27:72]
  wire [55:0] _T_119 = rdataSel[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_120 = {_T_119,rdataSel[7:0]}; // @[Cat.scala 30:58]
  wire [47:0] _T_124 = rdataSel[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_125 = {_T_124,rdataSel[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_129 = rdataSel[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_130 = {_T_129,rdataSel[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_132 = {56'h0,rdataSel[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_134 = {48'h0,rdataSel[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_136 = {32'h0,rdataSel[31:0]}; // @[Cat.scala 30:58]
  wire  _T_137 = 7'h0 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_138 = 7'h1 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_139 = 7'h2 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_140 = 7'h4 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_141 = 7'h5 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_142 = 7'h6 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_143 = _T_137 ? _T_120 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_144 = _T_138 ? _T_125 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_145 = _T_139 ? _T_130 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_146 = _T_140 ? _T_132 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_147 = _T_141 ? _T_134 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_148 = _T_142 ? _T_136 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_149 = _T_143 | _T_144; // @[Mux.scala 27:72]
  wire [63:0] _T_150 = _T_149 | _T_145; // @[Mux.scala 27:72]
  wire [63:0] _T_151 = _T_150 | _T_146; // @[Mux.scala 27:72]
  wire [63:0] _T_152 = _T_151 | _T_147; // @[Mux.scala 27:72]
  wire [63:0] rdataPartialLoad = _T_152 | _T_148; // @[Mux.scala 27:72]
  wire  _T_156 = ~io__in_bits_src1[0]; // @[UnpipelinedLSU.scala 416:27]
  wire  _T_158 = io__in_bits_src1[1:0] == 2'h0; // @[UnpipelinedLSU.scala 417:29]
  wire  _T_160 = io__in_bits_src1[2:0] == 3'h0; // @[UnpipelinedLSU.scala 418:29]
  wire  addrAligned = _T_26 | _T_27 & _T_156 | _T_28 & _T_158 | _T_29 & _T_160; // @[Mux.scala 27:72]
  wire  _T_178 = ~addrAligned; // @[UnpipelinedLSU.scala 429:60]
  wire  _T_196 = ~io__dmem_req_bits_cmd[0] & ~io__dmem_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_197 = io__dmem_req_valid & _T_196; // @[SimpleBus.scala 104:29]
  wire  _T_199 = _T_197 & _T_4; // @[UnpipelinedLSU.scala 434:39]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_9 = _T_197 | REG_1; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_208 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_11 = _T_208 | REG_2; // @[StopWatch.scala 24:20 30:{20,24}]
  assign io__out_valid = DTLBPF & state != 2'h0 | io__loadAddrMisaligned | io__storeAddrMisaligned | _T_64; // @[UnpipelinedLSU.scala 382:22]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 421:21]
  assign io__dmem_req_valid = io__in_valid & state == 2'h0 & ~io__loadAddrMisaligned & ~io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 379:75]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[UnpipelinedLSU.scala 370:68]
  assign io__dmem_req_bits_size = {{1'd0}, size}; // @[SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _T_35 | _T_33; // @[Mux.scala 27:72]
  assign io__dmem_resp_ready = 1'h1; // @[UnpipelinedLSU.scala 380:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF; // @[UnpipelinedLSU.scala 349:13]
  assign io__loadAddrMisaligned = io__in_valid & _T_1 & ~ISAMO2 & ~addrAligned; // @[UnpipelinedLSU.scala 429:57]
  assign io__storeAddrMisaligned = io__in_valid & (isStore | ISAMO2) & _T_178; // @[UnpipelinedLSU.scala 430:57]
  assign io_in_bits_src1 = io__in_bits_src1;
  always @(posedge clock) begin
    addrLatch <= io__in_bits_src1; // @[UnpipelinedLSU.scala 333:26]
    if (reset) begin // @[UnpipelinedLSU.scala 338:22]
      state <= 2'h0; // @[UnpipelinedLSU.scala 338:22]
    end else if (2'h0 == state) begin // @[UnpipelinedLSU.scala 351:18]
      if (_T_4 & ~DTLBENABLE) begin // @[UnpipelinedLSU.scala 354:45]
        state <= 2'h2; // @[UnpipelinedLSU.scala 354:53]
      end else if (_T_4 & DTLBENABLE) begin // @[UnpipelinedLSU.scala 353:45]
        state <= 2'h1; // @[UnpipelinedLSU.scala 353:53]
      end
    end else if (2'h1 == state) begin // @[UnpipelinedLSU.scala 351:18]
      if (DTLBFINISH & ~DTLBPF) begin // @[UnpipelinedLSU.scala 359:36]
        state <= 2'h2; // @[UnpipelinedLSU.scala 359:44]
      end else begin
        state <= _GEN_2;
      end
    end else if (2'h2 == state) begin // @[UnpipelinedLSU.scala 351:18]
      state <= _GEN_4;
    end else begin
      state <= _GEN_5;
    end
    rdataLatch <= io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 388:27]
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_14) begin // @[StopWatch.scala 31:19]
      REG_1 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_1 <= _GEN_9;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_14) begin // @[StopWatch.scala 31:19]
      REG_2 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_2 <= _GEN_11;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addrLatch = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  rdataLatch = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AtomALU(
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [6:0]  io_func,
  input         io_isWordOp,
  output [63:0] io_result
);
  wire  isAdderSub = ~io_func[6]; // @[LSU.scala 184:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_src2 ^ _T_2; // @[LSU.scala 185:33]
  wire [64:0] _T_4 = io_src1 + _T_3; // @[LSU.scala 185:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[LSU.scala 185:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[LSU.scala 185:60]
  wire [63:0] xorRes = io_src1 ^ io_src2; // @[LSU.scala 186:21]
  wire  sltu = ~adderRes[64]; // @[LSU.scala 187:14]
  wire  slt = xorRes[63] ^ sltu; // @[LSU.scala 188:28]
  wire [63:0] _T_9 = io_src1 & io_src2; // @[LSU.scala 194:32]
  wire [63:0] _T_10 = io_src1 | io_src2; // @[LSU.scala 195:32]
  wire [63:0] _T_12 = slt ? io_src1 : io_src2; // @[LSU.scala 196:29]
  wire [63:0] _T_14 = slt ? io_src2 : io_src1; // @[LSU.scala 197:29]
  wire [63:0] _T_16 = sltu ? io_src1 : io_src2; // @[LSU.scala 198:29]
  wire [63:0] _T_18 = sltu ? io_src2 : io_src1; // @[LSU.scala 199:29]
  wire [64:0] _T_20 = 6'h22 == io_func[5:0] ? {{1'd0}, io_src2} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_22 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _T_20; // @[Mux.scala 80:57]
  wire [64:0] _T_24 = 6'h25 == io_func[5:0] ? {{1'd0}, _T_9} : _T_22; // @[Mux.scala 80:57]
  wire [64:0] _T_26 = 6'h26 == io_func[5:0] ? {{1'd0}, _T_10} : _T_24; // @[Mux.scala 80:57]
  wire [64:0] _T_28 = 6'h37 == io_func[5:0] ? {{1'd0}, _T_12} : _T_26; // @[Mux.scala 80:57]
  wire [64:0] _T_30 = 6'h30 == io_func[5:0] ? {{1'd0}, _T_14} : _T_28; // @[Mux.scala 80:57]
  wire [64:0] _T_32 = 6'h31 == io_func[5:0] ? {{1'd0}, _T_16} : _T_30; // @[Mux.scala 80:57]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _T_18} : _T_32; // @[Mux.scala 80:57]
  wire [31:0] _T_37 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_38 = {_T_37,res[31:0]}; // @[Cat.scala 30:58]
  assign io_result = io_isWordOp ? _T_38 : res[63:0]; // @[LSU.scala 202:20]
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [63:0] io__in_bits_src2,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__wdata,
  input  [31:0] io__instr,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  output        setLr_0,
  input         DTLBPF,
  output        amoReq_0,
  input         DTLBENABLE,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH,
  output [63:0] setLrAddr_0,
  output        setLrVal_0,
  input  [63:0] lr_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_reset; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__in_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[UnpipelinedLSU.scala 47:28]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__wdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 47:28]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 47:28]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 47:28]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__isMMIO; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBPF; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBENABLE; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_ISAMO2; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io_in_bits_src1; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBFINISH; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] atomALU_io_src1; // @[UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_src2; // @[UnpipelinedLSU.scala 98:25]
  wire [6:0] atomALU_io_func; // @[UnpipelinedLSU.scala 98:25]
  wire  atomALU_io_isWordOp; // @[UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_result; // @[UnpipelinedLSU.scala 98:25]
  wire  atomReq = io__in_valid & io__in_bits_func[5]; // @[UnpipelinedLSU.scala 53:26]
  wire  _T_8 = io__in_bits_func == 7'h20; // @[LSU.scala 57:37]
  wire  _T_11 = io__in_bits_func == 7'h21; // @[LSU.scala 58:37]
  wire  _T_13 = io__in_bits_func[5] & ~_T_8 & ~_T_11; // @[LSU.scala 59:61]
  wire  amoReq = io__in_valid & _T_13; // @[UnpipelinedLSU.scala 54:26]
  wire  lrReq = io__in_valid & _T_8; // @[UnpipelinedLSU.scala 55:25]
  wire  scReq = io__in_valid & _T_11; // @[UnpipelinedLSU.scala 56:25]
  wire [2:0] funct3 = io__instr[14:12]; // @[UnpipelinedLSU.scala 64:26]
  wire  scInvalid = ~(io__in_bits_src1 == lr_addr) & scReq; // @[UnpipelinedLSU.scala 81:40]
  reg [2:0] state; // @[UnpipelinedLSU.scala 95:24]
  reg [63:0] atomMemReg; // @[UnpipelinedLSU.scala 96:25]
  reg [63:0] atomRegReg; // @[UnpipelinedLSU.scala 97:25]
  wire  _T_19 = 3'h0 == state; // @[UnpipelinedLSU.scala 128:20]
  wire  _T_22 = ~atomReq; // @[UnpipelinedLSU.scala 141:56]
  wire [63:0] _T_25 = io__in_bits_src1 + io__in_bits_src2; // @[UnpipelinedLSU.scala 143:46]
  wire  _T_26 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_1 = amoReq ? 3'h5 : 3'h0; // @[UnpipelinedLSU.scala 149:17 152:{21,28}]
  wire [2:0] _GEN_2 = lrReq ? 3'h3 : _GEN_1; // @[UnpipelinedLSU.scala 153:{20,27}]
  wire [2:0] _T_29 = scInvalid ? 3'h0 : 3'h4; // @[UnpipelinedLSU.scala 154:33]
  wire  _T_30 = 3'h1 == state; // @[UnpipelinedLSU.scala 128:20]
  wire [2:0] _GEN_4 = io__out_valid ? 3'h0 : state; // @[UnpipelinedLSU.scala 168:{28,35} 95:24]
  wire [1:0] _T_44 = funct3[0] ? 2'h3 : 2'h2; // @[UnpipelinedLSU.scala 188:42]
  wire [2:0] _GEN_5 = _T_26 ? 3'h6 : state; // @[UnpipelinedLSU.scala 192:39 193:17 95:24]
  wire [3:0] _T_48 = funct3[0] ? 4'hb : 4'ha; // @[UnpipelinedLSU.scala 219:42]
  wire [2:0] _GEN_6 = _T_26 ? 3'h0 : state; // @[UnpipelinedLSU.scala 223:39 224:17 95:24]
  wire [63:0] _GEN_11 = io__in_bits_src1; // @[UnpipelinedLSU.scala 128:20 245:36]
  wire  _GEN_14 = 3'h4 == state & _T_26; // @[UnpipelinedLSU.scala 128:20 126:32 249:36]
  wire [2:0] _GEN_16 = 3'h4 == state ? _GEN_6 : state; // @[UnpipelinedLSU.scala 128:20 95:24]
  wire  _GEN_17 = 3'h3 == state | 3'h4 == state; // @[UnpipelinedLSU.scala 128:20 229:36]
  wire [3:0] _GEN_20 = 3'h3 == state ? {{2'd0}, _T_44} : _T_48; // @[UnpipelinedLSU.scala 128:20 233:36]
  wire  _GEN_22 = 3'h3 == state ? _T_26 : _GEN_14; // @[UnpipelinedLSU.scala 128:20 235:36]
  wire [2:0] _GEN_24 = 3'h3 == state ? _GEN_6 : _GEN_16; // @[UnpipelinedLSU.scala 128:20]
  wire  _GEN_25 = 3'h7 == state | _GEN_17; // @[UnpipelinedLSU.scala 128:20 215:36]
  wire [3:0] _GEN_28 = 3'h7 == state ? _T_48 : _GEN_20; // @[UnpipelinedLSU.scala 128:20 219:36]
  wire [63:0] _GEN_29 = 3'h7 == state ? atomMemReg : io__wdata; // @[UnpipelinedLSU.scala 128:20 220:36]
  wire  _GEN_30 = 3'h7 == state ? _T_26 : _GEN_22; // @[UnpipelinedLSU.scala 128:20 221:36]
  wire [2:0] _GEN_32 = 3'h7 == state ? _GEN_6 : _GEN_24; // @[UnpipelinedLSU.scala 128:20]
  wire  _GEN_33 = 3'h6 == state ? 1'h0 : _GEN_25; // @[UnpipelinedLSU.scala 128:20 201:36]
  wire  _GEN_34 = 3'h6 == state ? 1'h0 : 1'h1; // @[UnpipelinedLSU.scala 128:20 202:36]
  wire  _GEN_38 = 3'h6 == state ? 1'h0 : _GEN_30; // @[UnpipelinedLSU.scala 128:20 207:36]
  wire [2:0] _GEN_40 = 3'h6 == state ? 3'h7 : _GEN_32; // @[UnpipelinedLSU.scala 128:20 209:15]
  wire  _GEN_42 = 3'h5 == state | _GEN_33; // @[UnpipelinedLSU.scala 128:20 184:36]
  wire  _GEN_43 = 3'h5 == state | _GEN_34; // @[UnpipelinedLSU.scala 128:20 185:36]
  wire [3:0] _GEN_45 = 3'h5 == state ? {{2'd0}, _T_44} : _GEN_28; // @[UnpipelinedLSU.scala 128:20 188:36]
  wire  _GEN_47 = 3'h5 == state ? 1'h0 : _GEN_38; // @[UnpipelinedLSU.scala 128:20 190:36]
  wire [2:0] _GEN_49 = 3'h5 == state ? _GEN_5 : _GEN_40; // @[UnpipelinedLSU.scala 128:20]
  wire  _GEN_52 = 3'h1 == state | _GEN_42; // @[UnpipelinedLSU.scala 128:20 159:36]
  wire  _GEN_53 = 3'h1 == state | _GEN_43; // @[UnpipelinedLSU.scala 128:20 160:36]
  wire [6:0] _GEN_55 = 3'h1 == state ? io__in_bits_func : {{3'd0}, _GEN_45}; // @[UnpipelinedLSU.scala 128:20 163:36]
  wire [63:0] _GEN_56 = 3'h1 == state ? io__wdata : _GEN_29; // @[UnpipelinedLSU.scala 128:20 164:36]
  wire  _GEN_58 = 3'h1 == state ? lsExecUnit_io__out_valid : _GEN_47; // @[UnpipelinedLSU.scala 128:20 166:36]
  wire  _GEN_68 = 3'h0 == state ? lsExecUnit_io__out_valid | scInvalid : _GEN_58; // @[UnpipelinedLSU.scala 128:20 148:38]
  wire [63:0] _T_68 = state == 3'h7 ? atomRegReg : lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 275:45]
  wire  setLr = io__out_valid & (lrReq | scReq); // @[UnpipelinedLSU.scala 270:28]
  wire  setLrVal = lrReq; // @[UnpipelinedLSU.scala 55:25]
  wire [63:0] setLrAddr = io__in_bits_src1; // @[UnpipelinedLSU.scala 272:15 72:25]
  LSExecUnit lsExecUnit ( // @[UnpipelinedLSU.scala 47:28]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__loadAddrMisaligned(lsExecUnit_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsExecUnit_io__storeAddrMisaligned),
    .DTLBPF(lsExecUnit_DTLBPF),
    .DTLBENABLE(lsExecUnit_DTLBENABLE),
    .ISAMO2(lsExecUnit_ISAMO2),
    .io_in_bits_src1(lsExecUnit_io_in_bits_src1),
    .DTLBFINISH(lsExecUnit_DTLBFINISH)
  );
  AtomALU atomALU ( // @[UnpipelinedLSU.scala 98:25]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io__out_valid = DTLBPF | io__loadAddrMisaligned | io__storeAddrMisaligned | _GEN_68; // @[UnpipelinedLSU.scala 257:68 259:20]
  assign io__out_bits = scReq ? {{63'd0}, scInvalid} : _T_68; // @[UnpipelinedLSU.scala 275:23]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 274:13]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 49:15]
  assign io__loadAddrMisaligned = lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 285:27]
  assign io__storeAddrMisaligned = lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 286:28]
  assign setLr_0 = setLr;
  assign amoReq_0 = amoReq;
  assign io_in_bits_src1 = lsExecUnit_io_in_bits_src1;
  assign setLrAddr_0 = _GEN_11;
  assign setLrVal_0 = setLrVal;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = 3'h0 == state ? io__in_valid & ~atomReq : _GEN_52; // @[UnpipelinedLSU.scala 128:20 141:38]
  assign lsExecUnit_io__in_bits_src1 = 3'h0 == state ? _T_25 : io__in_bits_src1; // @[UnpipelinedLSU.scala 128:20 143:38]
  assign lsExecUnit_io__in_bits_func = 3'h0 == state ? io__in_bits_func : _GEN_55; // @[UnpipelinedLSU.scala 128:20 145:38]
  assign lsExecUnit_io__out_ready = 3'h0 == state | _GEN_53; // @[UnpipelinedLSU.scala 128:20 142:38]
  assign lsExecUnit_io__wdata = 3'h0 == state ? io__wdata : _GEN_56; // @[UnpipelinedLSU.scala 128:20 146:38]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_DTLBPF = DTLBPF;
  assign lsExecUnit_DTLBENABLE = DTLBENABLE;
  assign lsExecUnit_ISAMO2 = amoReq;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign atomALU_io_src1 = atomMemReg; // @[UnpipelinedLSU.scala 99:21]
  assign atomALU_io_src2 = io__wdata; // @[UnpipelinedLSU.scala 100:21]
  assign atomALU_io_func = io__in_bits_func; // @[UnpipelinedLSU.scala 101:21]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[UnpipelinedLSU.scala 66:22]
  always @(posedge clock) begin
    if (reset) begin // @[UnpipelinedLSU.scala 95:24]
      state <= 3'h0; // @[UnpipelinedLSU.scala 95:24]
    end else if (DTLBPF | io__loadAddrMisaligned | io__storeAddrMisaligned) begin // @[UnpipelinedLSU.scala 257:68]
      state <= 3'h0; // @[UnpipelinedLSU.scala 258:13]
    end else if (3'h0 == state) begin // @[UnpipelinedLSU.scala 128:20]
      if (scReq) begin // @[UnpipelinedLSU.scala 154:20]
        state <= _T_29; // @[UnpipelinedLSU.scala 154:27]
      end else begin
        state <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[UnpipelinedLSU.scala 128:20]
      state <= _GEN_4;
    end else begin
      state <= _GEN_49;
    end
    if (!(3'h0 == state)) begin // @[UnpipelinedLSU.scala 128:20]
      if (!(3'h1 == state)) begin // @[UnpipelinedLSU.scala 128:20]
        if (3'h5 == state) begin // @[UnpipelinedLSU.scala 128:20]
          atomMemReg <= lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 196:20]
        end else if (3'h6 == state) begin // @[UnpipelinedLSU.scala 128:20]
          atomMemReg <= atomALU_io_result; // @[UnpipelinedLSU.scala 210:20]
        end
      end
    end
    if (!(3'h0 == state)) begin // @[UnpipelinedLSU.scala 128:20]
      if (!(3'h1 == state)) begin // @[UnpipelinedLSU.scala 128:20]
        if (3'h5 == state) begin // @[UnpipelinedLSU.scala 128:20]
          atomRegReg <= lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 197:20]
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_19 & _T_30 & ~(_T_22 | ~amoReq | ~lrReq | ~scReq | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UnpipelinedLSU.scala:167 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[UnpipelinedLSU.scala 167:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_19 & _T_30 & ~(_T_22 | ~amoReq | ~lrReq | ~scReq | reset)) begin
          $fatal; // @[UnpipelinedLSU.scala 167:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  atomMemReg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  atomRegReg = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [64:0]  io_in_bits_0,
  input  [64:0]  io_in_bits_1,
  input          io_out_ready,
  output         io_out_valid,
  output [129:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] REG; // @[MDU.scala 56:43]
  reg [64:0] REG_1; // @[MDU.scala 56:43]
  reg [129:0] REG_2; // @[MDU.scala 57:60]
  reg [129:0] REG_3; // @[MDU.scala 57:52]
  reg [129:0] REG_4; // @[MDU.scala 57:44]
  reg  REG_5; // @[MDU.scala 56:43]
  reg  REG_6; // @[MDU.scala 57:60]
  reg  REG_7; // @[MDU.scala 57:52]
  reg  REG_8; // @[MDU.scala 57:44]
  reg  busy; // @[MDU.scala 62:21]
  wire  _GEN_0 = io_in_valid & ~busy | busy; // @[MDU.scala 62:21 63:{31,38}]
  assign io_in_ready = ~busy; // @[MDU.scala 65:49]
  assign io_out_valid = REG_8; // @[MDU.scala 60:16]
  assign io_out_bits = REG_4; // @[MDU.scala 59:37]
  always @(posedge clock) begin
    REG <= io_in_bits_0; // @[MDU.scala 56:43]
    REG_1 <= io_in_bits_1; // @[MDU.scala 56:43]
    REG_2 <= $signed(REG) * $signed(REG_1); // @[MDU.scala 58:49]
    REG_3 <= REG_2; // @[MDU.scala 57:52]
    REG_4 <= REG_3; // @[MDU.scala 57:44]
    REG_5 <= io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
    REG_6 <= REG_5; // @[MDU.scala 57:60]
    REG_7 <= REG_6; // @[MDU.scala 57:52]
    REG_8 <= REG_7; // @[MDU.scala 57:44]
    if (reset) begin // @[MDU.scala 62:21]
      busy <= 1'h0; // @[MDU.scala 62:21]
    end else if (io_out_valid) begin // @[MDU.scala 64:23]
      busy <= 1'h0; // @[MDU.scala 64:30]
    end else begin
      busy <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  REG = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  REG_1 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  REG_2 = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  REG_3 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  REG_4 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  REG_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [63:0]  io_in_bits_0,
  input  [63:0]  io_in_bits_1,
  input          io_sign,
  output         io_out_valid,
  output [127:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[MDU.scala 77:22]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  newReq = state == 3'h0 & _T_1; // @[MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[MDU.scala 81:18]
  reg [128:0] shiftReg; // @[MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[MDU.scala 72:24]
  wire [63:0] _T_4 = 64'h0 - io_in_bits_0; // @[MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_4 : io_in_bits_0; // @[MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[MDU.scala 72:24]
  wire [63:0] _T_7 = 64'h0 - io_in_bits_1; // @[MDU.scala 73:16]
  reg  aSignReg; // @[Reg.scala 15:16]
  wire  _T_10 = (aSign ^ bSign) & ~divBy0; // @[MDU.scala 90:44]
  reg  qSignReg; // @[Reg.scala 15:16]
  reg [63:0] bReg; // @[Reg.scala 15:16]
  wire [64:0] _T_11 = {aVal,1'h0}; // @[Cat.scala 30:58]
  reg [64:0] aValx2Reg; // @[Reg.scala 15:16]
  reg [5:0] value; // @[Counter.scala 60:40]
  wire [31:0] hi_1 = bReg[63:32]; // @[CircuitMath.scala 35:17]
  wire [31:0] lo_1 = bReg[31:0]; // @[CircuitMath.scala 36:17]
  wire  useHi = |hi_1; // @[CircuitMath.scala 37:22]
  wire [15:0] hi_2 = hi_1[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_2 = hi_1[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_1 = |hi_2; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_3 = hi_2[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_3 = hi_2[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_2 = |hi_3; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_4 = hi_3[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_4 = hi_3[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_3 = |hi_4; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_16 = hi_4[2] ? 2'h2 : {{1'd0}, hi_4[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_17 = hi_4[3] ? 2'h3 : _T_16; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_21 = lo_4[2] ? 2'h2 : {{1'd0}, lo_4[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_22 = lo_4[3] ? 2'h3 : _T_21; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_23 = useHi_3 ? _T_17 : _T_22; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_24 = {useHi_3,_T_23}; // @[Cat.scala 30:58]
  wire [3:0] hi_5 = lo_3[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_5 = lo_3[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_4 = |hi_5; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_28 = hi_5[2] ? 2'h2 : {{1'd0}, hi_5[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_29 = hi_5[3] ? 2'h3 : _T_28; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_33 = lo_5[2] ? 2'h2 : {{1'd0}, lo_5[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_34 = lo_5[3] ? 2'h3 : _T_33; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_35 = useHi_4 ? _T_29 : _T_34; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_36 = {useHi_4,_T_35}; // @[Cat.scala 30:58]
  wire [2:0] _T_37 = useHi_2 ? _T_24 : _T_36; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_38 = {useHi_2,_T_37}; // @[Cat.scala 30:58]
  wire [7:0] hi_6 = lo_2[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_6 = lo_2[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_5 = |hi_6; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_7 = hi_6[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_7 = hi_6[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_6 = |hi_7; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_42 = hi_7[2] ? 2'h2 : {{1'd0}, hi_7[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_43 = hi_7[3] ? 2'h3 : _T_42; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_47 = lo_7[2] ? 2'h2 : {{1'd0}, lo_7[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_48 = lo_7[3] ? 2'h3 : _T_47; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_49 = useHi_6 ? _T_43 : _T_48; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_50 = {useHi_6,_T_49}; // @[Cat.scala 30:58]
  wire [3:0] hi_8 = lo_6[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_8 = lo_6[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_7 = |hi_8; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_54 = hi_8[2] ? 2'h2 : {{1'd0}, hi_8[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_55 = hi_8[3] ? 2'h3 : _T_54; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_59 = lo_8[2] ? 2'h2 : {{1'd0}, lo_8[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_60 = lo_8[3] ? 2'h3 : _T_59; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_61 = useHi_7 ? _T_55 : _T_60; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_62 = {useHi_7,_T_61}; // @[Cat.scala 30:58]
  wire [2:0] _T_63 = useHi_5 ? _T_50 : _T_62; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_64 = {useHi_5,_T_63}; // @[Cat.scala 30:58]
  wire [3:0] _T_65 = useHi_1 ? _T_38 : _T_64; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_66 = {useHi_1,_T_65}; // @[Cat.scala 30:58]
  wire [15:0] hi_9 = lo_1[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_9 = lo_1[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_8 = |hi_9; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_10 = hi_9[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_10 = hi_9[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_9 = |hi_10; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_11 = hi_10[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_11 = hi_10[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_10 = |hi_11; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_70 = hi_11[2] ? 2'h2 : {{1'd0}, hi_11[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_71 = hi_11[3] ? 2'h3 : _T_70; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_75 = lo_11[2] ? 2'h2 : {{1'd0}, lo_11[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_76 = lo_11[3] ? 2'h3 : _T_75; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_77 = useHi_10 ? _T_71 : _T_76; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_78 = {useHi_10,_T_77}; // @[Cat.scala 30:58]
  wire [3:0] hi_12 = lo_10[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_12 = lo_10[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_11 = |hi_12; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_82 = hi_12[2] ? 2'h2 : {{1'd0}, hi_12[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_83 = hi_12[3] ? 2'h3 : _T_82; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_87 = lo_12[2] ? 2'h2 : {{1'd0}, lo_12[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_88 = lo_12[3] ? 2'h3 : _T_87; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_89 = useHi_11 ? _T_83 : _T_88; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_90 = {useHi_11,_T_89}; // @[Cat.scala 30:58]
  wire [2:0] _T_91 = useHi_9 ? _T_78 : _T_90; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_92 = {useHi_9,_T_91}; // @[Cat.scala 30:58]
  wire [7:0] hi_13 = lo_9[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_13 = lo_9[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_12 = |hi_13; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_14 = hi_13[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_14 = hi_13[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_13 = |hi_14; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_96 = hi_14[2] ? 2'h2 : {{1'd0}, hi_14[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_97 = hi_14[3] ? 2'h3 : _T_96; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_101 = lo_14[2] ? 2'h2 : {{1'd0}, lo_14[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_102 = lo_14[3] ? 2'h3 : _T_101; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_103 = useHi_13 ? _T_97 : _T_102; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_104 = {useHi_13,_T_103}; // @[Cat.scala 30:58]
  wire [3:0] hi_15 = lo_13[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_15 = lo_13[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_14 = |hi_15; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_108 = hi_15[2] ? 2'h2 : {{1'd0}, hi_15[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_109 = hi_15[3] ? 2'h3 : _T_108; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_113 = lo_15[2] ? 2'h2 : {{1'd0}, lo_15[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_114 = lo_15[3] ? 2'h3 : _T_113; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_115 = useHi_14 ? _T_109 : _T_114; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_116 = {useHi_14,_T_115}; // @[Cat.scala 30:58]
  wire [2:0] _T_117 = useHi_12 ? _T_104 : _T_116; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_118 = {useHi_12,_T_117}; // @[Cat.scala 30:58]
  wire [3:0] _T_119 = useHi_8 ? _T_92 : _T_118; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_120 = {useHi_8,_T_119}; // @[Cat.scala 30:58]
  wire [4:0] _T_121 = useHi ? _T_66 : _T_120; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_122 = {useHi,_T_121}; // @[Cat.scala 30:58]
  wire [6:0] _GEN_18 = {{1'd0}, _T_122}; // @[MDU.scala 105:31]
  wire [6:0] _T_123 = 7'h40 | _GEN_18; // @[MDU.scala 105:31]
  wire  hi_16 = aValx2Reg[64]; // @[CircuitMath.scala 35:17]
  wire [63:0] lo_16 = aValx2Reg[63:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_15 = |hi_16; // @[CircuitMath.scala 37:22]
  wire [31:0] hi_17 = lo_16[63:32]; // @[CircuitMath.scala 35:17]
  wire [31:0] lo_17 = lo_16[31:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_16 = |hi_17; // @[CircuitMath.scala 37:22]
  wire [15:0] hi_18 = hi_17[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_18 = hi_17[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_17 = |hi_18; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_19 = hi_18[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_19 = hi_18[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_18 = |hi_19; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_20 = hi_19[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_20 = hi_19[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_19 = |hi_20; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_127 = hi_20[2] ? 2'h2 : {{1'd0}, hi_20[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_128 = hi_20[3] ? 2'h3 : _T_127; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_132 = lo_20[2] ? 2'h2 : {{1'd0}, lo_20[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_133 = lo_20[3] ? 2'h3 : _T_132; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_134 = useHi_19 ? _T_128 : _T_133; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_135 = {useHi_19,_T_134}; // @[Cat.scala 30:58]
  wire [3:0] hi_21 = lo_19[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_21 = lo_19[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_20 = |hi_21; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_139 = hi_21[2] ? 2'h2 : {{1'd0}, hi_21[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_140 = hi_21[3] ? 2'h3 : _T_139; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_144 = lo_21[2] ? 2'h2 : {{1'd0}, lo_21[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_145 = lo_21[3] ? 2'h3 : _T_144; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_146 = useHi_20 ? _T_140 : _T_145; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_147 = {useHi_20,_T_146}; // @[Cat.scala 30:58]
  wire [2:0] _T_148 = useHi_18 ? _T_135 : _T_147; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_149 = {useHi_18,_T_148}; // @[Cat.scala 30:58]
  wire [7:0] hi_22 = lo_18[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_22 = lo_18[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_21 = |hi_22; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_23 = hi_22[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_23 = hi_22[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_22 = |hi_23; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_153 = hi_23[2] ? 2'h2 : {{1'd0}, hi_23[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_154 = hi_23[3] ? 2'h3 : _T_153; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_158 = lo_23[2] ? 2'h2 : {{1'd0}, lo_23[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_159 = lo_23[3] ? 2'h3 : _T_158; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_160 = useHi_22 ? _T_154 : _T_159; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_161 = {useHi_22,_T_160}; // @[Cat.scala 30:58]
  wire [3:0] hi_24 = lo_22[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_24 = lo_22[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_23 = |hi_24; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_165 = hi_24[2] ? 2'h2 : {{1'd0}, hi_24[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_166 = hi_24[3] ? 2'h3 : _T_165; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_170 = lo_24[2] ? 2'h2 : {{1'd0}, lo_24[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_171 = lo_24[3] ? 2'h3 : _T_170; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_172 = useHi_23 ? _T_166 : _T_171; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_173 = {useHi_23,_T_172}; // @[Cat.scala 30:58]
  wire [2:0] _T_174 = useHi_21 ? _T_161 : _T_173; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_175 = {useHi_21,_T_174}; // @[Cat.scala 30:58]
  wire [3:0] _T_176 = useHi_17 ? _T_149 : _T_175; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_177 = {useHi_17,_T_176}; // @[Cat.scala 30:58]
  wire [15:0] hi_25 = lo_17[31:16]; // @[CircuitMath.scala 35:17]
  wire [15:0] lo_25 = lo_17[15:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_24 = |hi_25; // @[CircuitMath.scala 37:22]
  wire [7:0] hi_26 = hi_25[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_26 = hi_25[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_25 = |hi_26; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_27 = hi_26[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_27 = hi_26[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_26 = |hi_27; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_181 = hi_27[2] ? 2'h2 : {{1'd0}, hi_27[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_182 = hi_27[3] ? 2'h3 : _T_181; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_186 = lo_27[2] ? 2'h2 : {{1'd0}, lo_27[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_187 = lo_27[3] ? 2'h3 : _T_186; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_188 = useHi_26 ? _T_182 : _T_187; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_189 = {useHi_26,_T_188}; // @[Cat.scala 30:58]
  wire [3:0] hi_28 = lo_26[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_28 = lo_26[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_27 = |hi_28; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_193 = hi_28[2] ? 2'h2 : {{1'd0}, hi_28[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_194 = hi_28[3] ? 2'h3 : _T_193; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_198 = lo_28[2] ? 2'h2 : {{1'd0}, lo_28[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_199 = lo_28[3] ? 2'h3 : _T_198; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_200 = useHi_27 ? _T_194 : _T_199; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_201 = {useHi_27,_T_200}; // @[Cat.scala 30:58]
  wire [2:0] _T_202 = useHi_25 ? _T_189 : _T_201; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_203 = {useHi_25,_T_202}; // @[Cat.scala 30:58]
  wire [7:0] hi_29 = lo_25[15:8]; // @[CircuitMath.scala 35:17]
  wire [7:0] lo_29 = lo_25[7:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_28 = |hi_29; // @[CircuitMath.scala 37:22]
  wire [3:0] hi_30 = hi_29[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_30 = hi_29[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_29 = |hi_30; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_207 = hi_30[2] ? 2'h2 : {{1'd0}, hi_30[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_208 = hi_30[3] ? 2'h3 : _T_207; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_212 = lo_30[2] ? 2'h2 : {{1'd0}, lo_30[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_213 = lo_30[3] ? 2'h3 : _T_212; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_214 = useHi_29 ? _T_208 : _T_213; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_215 = {useHi_29,_T_214}; // @[Cat.scala 30:58]
  wire [3:0] hi_31 = lo_29[7:4]; // @[CircuitMath.scala 35:17]
  wire [3:0] lo_31 = lo_29[3:0]; // @[CircuitMath.scala 36:17]
  wire  useHi_30 = |hi_31; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_219 = hi_31[2] ? 2'h2 : {{1'd0}, hi_31[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_220 = hi_31[3] ? 2'h3 : _T_219; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_224 = lo_31[2] ? 2'h2 : {{1'd0}, lo_31[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_225 = lo_31[3] ? 2'h3 : _T_224; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_226 = useHi_30 ? _T_220 : _T_225; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_227 = {useHi_30,_T_226}; // @[Cat.scala 30:58]
  wire [2:0] _T_228 = useHi_28 ? _T_215 : _T_227; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_229 = {useHi_28,_T_228}; // @[Cat.scala 30:58]
  wire [3:0] _T_230 = useHi_24 ? _T_203 : _T_229; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_231 = {useHi_24,_T_230}; // @[Cat.scala 30:58]
  wire [4:0] _T_232 = useHi_16 ? _T_177 : _T_231; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_233 = {useHi_16,_T_232}; // @[Cat.scala 30:58]
  wire [5:0] _T_234 = useHi_15 ? 6'h0 : _T_233; // @[CircuitMath.scala 38:21]
  wire [6:0] _T_235 = {useHi_15,_T_234}; // @[Cat.scala 30:58]
  wire [6:0] _T_237 = _T_123 - _T_235; // @[MDU.scala 105:45]
  wire [6:0] _value_T_1 = _T_237 >= 7'h3f ? 7'h3f : _T_237; // @[MDU.scala 109:38]
  wire [6:0] _value_T_2 = divBy0 ? 7'h0 : _value_T_1; // @[MDU.scala 109:21]
  wire [127:0] _GEN_0 = {{63'd0}, aValx2Reg}; // @[MDU.scala 112:27]
  wire [127:0] _T_239 = _GEN_0 << value; // @[MDU.scala 112:27]
  wire [64:0] _GEN_19 = {{1'd0}, bReg}; // @[MDU.scala 115:28]
  wire  _T_241 = hi >= _GEN_19; // @[MDU.scala 115:28]
  wire [64:0] _T_243 = hi - _GEN_19; // @[MDU.scala 116:36]
  wire [64:0] _T_244 = _T_241 ? _T_243 : hi; // @[MDU.scala 116:24]
  wire [128:0] _T_246 = {_T_244[63:0],lo,_T_241}; // @[Cat.scala 30:58]
  wire  wrap = value == 6'h3f; // @[Counter.scala 72:24]
  wire [5:0] _value_T_4 = value + 6'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_4 = wrap ? 3'h4 : state; // @[MDU.scala 118:{36,44} 77:22]
  wire [2:0] _GEN_5 = state == 3'h4 ? 3'h0 : state; // @[MDU.scala 119:36 120:11 77:22]
  wire [5:0] _GEN_7 = state == 3'h3 ? _value_T_4 : value; // @[MDU.scala 114:37 Counter.scala 76:15 60:40]
  wire [2:0] _GEN_8 = state == 3'h3 ? _GEN_4 : _GEN_5; // @[MDU.scala 114:37]
  wire [5:0] _GEN_11 = state == 3'h2 ? value : _GEN_7; // @[MDU.scala 111:35 Counter.scala 60:40]
  wire [6:0] _GEN_12 = state == 3'h1 ? _value_T_2 : {{1'd0}, _GEN_11}; // @[MDU.scala 109:15 97:34]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, value} : _GEN_12; // @[MDU.scala 95:17 Counter.scala 60:40]
  wire [63:0] r = hi[64:1]; // @[MDU.scala 123:13]
  wire [63:0] _T_250 = 64'h0 - lo; // @[MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _T_250 : lo; // @[MDU.scala 124:17]
  wire [63:0] _T_252 = 64'h0 - r; // @[MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _T_252 : r; // @[MDU.scala 125:17]
  assign io_in_ready = state == 3'h0; // @[MDU.scala 129:25]
  assign io_out_valid = state == 3'h4; // @[MDU.scala 128:39]
  assign io_out_bits = {resR,resQ}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[MDU.scala 77:22]
      state <= 3'h0; // @[MDU.scala 77:22]
    end else if (newReq) begin // @[MDU.scala 95:17]
      state <= 3'h1; // @[MDU.scala 96:11]
    end else if (state == 3'h1) begin // @[MDU.scala 97:34]
      state <= 3'h2; // @[MDU.scala 110:11]
    end else if (state == 3'h2) begin // @[MDU.scala 111:35]
      state <= 3'h3; // @[MDU.scala 113:11]
    end else begin
      state <= _GEN_8;
    end
    if (!(newReq)) begin // @[MDU.scala 95:17]
      if (!(state == 3'h1)) begin // @[MDU.scala 97:34]
        if (state == 3'h2) begin // @[MDU.scala 111:35]
          shiftReg <= {{1'd0}, _T_239}; // @[MDU.scala 112:14]
        end else if (state == 3'h3) begin // @[MDU.scala 114:37]
          shiftReg <= _T_246; // @[MDU.scala 116:14]
        end
      end
    end
    if (newReq) begin // @[Reg.scala 16:19]
      aSignReg <= aSign; // @[Reg.scala 16:23]
    end
    if (newReq) begin // @[Reg.scala 16:19]
      qSignReg <= _T_10; // @[Reg.scala 16:23]
    end
    if (newReq) begin // @[Reg.scala 16:19]
      if (bSign) begin // @[MDU.scala 73:12]
        bReg <= _T_7;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin // @[Reg.scala 16:19]
      aValx2Reg <= _T_11; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 6'h0; // @[Counter.scala 60:40]
    end else begin
      value <= _GEN_16[5:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[MDU.scala 151:19]
  wire  mul_reset; // @[MDU.scala 151:19]
  wire  mul_io_in_ready; // @[MDU.scala 151:19]
  wire  mul_io_in_valid; // @[MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[MDU.scala 151:19]
  wire  mul_io_out_ready; // @[MDU.scala 151:19]
  wire  mul_io_out_valid; // @[MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[MDU.scala 151:19]
  wire  div_clock; // @[MDU.scala 152:19]
  wire  div_reset; // @[MDU.scala 152:19]
  wire  div_io_in_ready; // @[MDU.scala 152:19]
  wire  div_io_in_valid; // @[MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[MDU.scala 152:19]
  wire  div_io_sign; // @[MDU.scala 152:19]
  wire  div_io_out_valid; // @[MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[MDU.scala 43:25]
  wire [64:0] _T_4 = {1'h0,io_in_bits_src1}; // @[Cat.scala 30:58]
  wire [64:0] _T_6 = {io_in_bits_src1[63],io_in_bits_src1}; // @[Cat.scala 30:58]
  wire  _T_10 = 2'h0 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_11 = 2'h1 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_12 = 2'h2 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_13 = 2'h3 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [64:0] _T_14 = _T_10 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_15 = _T_11 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_16 = _T_12 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_17 = _T_13 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_18 = _T_14 | _T_15; // @[Mux.scala 27:72]
  wire [64:0] _T_19 = _T_18 | _T_16; // @[Mux.scala 27:72]
  wire [64:0] _T_22 = {1'h0,io_in_bits_src2}; // @[Cat.scala 30:58]
  wire [64:0] _T_24 = {io_in_bits_src2[63],io_in_bits_src2}; // @[Cat.scala 30:58]
  wire [64:0] _T_31 = _T_10 ? _T_22 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_32 = _T_11 ? _T_24 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_33 = _T_12 ? _T_22 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_34 = _T_13 ? _T_22 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_35 = _T_31 | _T_32; // @[Mux.scala 27:72]
  wire [64:0] _T_36 = _T_35 | _T_33; // @[Mux.scala 27:72]
  wire [31:0] _T_41 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_42 = {_T_41,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_44 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_45 = isDivSign ? _T_42 : _T_44; // @[MDU.scala 169:47]
  wire [31:0] _T_50 = io_in_bits_src2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_51 = {_T_50,io_in_bits_src2[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_53 = {32'h0,io_in_bits_src2[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_54 = isDivSign ? _T_51 : _T_53; // @[MDU.scala 169:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[MDU.scala 178:16]
  wire [31:0] _T_69 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_70 = {_T_69,res[31:0]}; // @[Cat.scala 30:58]
  wire  _T_72 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[MDU.scala 181:50]
  wire  isDivReg = _T_72 ? isDiv : REG; // @[MDU.scala 181:21]
  wire  _T_75 = mul_io_out_ready & mul_io_out_valid; // @[Decoupled.scala 40:37]
  Multiplier mul ( // @[MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[MDU.scala 182:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[MDU.scala 183:22]
  assign io_out_bits = isW ? _T_70 : res; // @[MDU.scala 179:21]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[MDU.scala 173:34]
  assign mul_io_in_bits_0 = _T_19 | _T_17; // @[Mux.scala 27:72]
  assign mul_io_in_bits_1 = _T_36 | _T_34; // @[Mux.scala 27:72]
  assign mul_io_out_ready = 1'h1; // @[MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[MDU.scala 174:34]
  assign div_io_in_bits_0 = isW ? _T_45 : io_in_bits_src1; // @[MDU.scala 169:38]
  assign div_io_in_bits_1 = isW ? _T_54 : io_in_bits_src2; // @[MDU.scala 169:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[MDU.scala 42:39]
  always @(posedge clock) begin
    REG <= io_in_bits_func[2]; // @[MDU.scala 41:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input         io_cfIn_exceptionVec_1,
  input         io_cfIn_exceptionVec_2,
  input         io_cfIn_exceptionVec_4,
  input         io_cfIn_exceptionVec_6,
  input         io_cfIn_exceptionVec_12,
  input         io_cfIn_intrVec_0,
  input         io_cfIn_intrVec_1,
  input         io_cfIn_intrVec_2,
  input         io_cfIn_intrVec_3,
  input         io_cfIn_intrVec_4,
  input         io_cfIn_intrVec_5,
  input         io_cfIn_intrVec_6,
  input         io_cfIn_intrVec_7,
  input         io_cfIn_intrVec_8,
  input         io_cfIn_intrVec_9,
  input         io_cfIn_intrVec_10,
  input         io_cfIn_intrVec_11,
  input         io_cfIn_crossPageIPFFix,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         io_instrValid,
  output [1:0]  io_imemMMU_priviledgeMode,
  output [1:0]  io_dmemMMU_priviledgeMode,
  output        io_dmemMMU_status_sum,
  output        io_dmemMMU_status_mxr,
  input         io_dmemMMU_loadPF,
  input         io_dmemMMU_storePF,
  input  [38:0] io_dmemMMU_addr,
  output        io_wenFix,
  input         set_lr,
  output [63:0] perfCnts_2_0,
  output [63:0] satp_0,
  input         perfCntCondMinstret,
  input         mtip_0,
  input         meip_0,
  input  [63:0] LSUADDR,
  output [11:0] intrVec_0,
  input         msip_0,
  input  [63:0] set_lr_addr,
  input         perfCntCondMultiCommit,
  input         set_lr_val,
  output [63:0] lrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtvec; // @[CSR.scala 252:22]
  reg [63:0] mcounteren; // @[CSR.scala 253:27]
  reg [63:0] mcause; // @[CSR.scala 254:23]
  reg [63:0] mtval; // @[CSR.scala 255:22]
  reg [63:0] mepc; // @[CSR.scala 256:17]
  reg [63:0] mie; // @[CSR.scala 258:20]
  reg [63:0] mipReg; // @[CSR.scala 260:24]
  wire [11:0] _T_1 = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[CSR.scala 262:22]
  wire [63:0] _GEN_78 = {{52'd0}, _T_1}; // @[CSR.scala 262:29]
  wire [63:0] _T_2 = _GEN_78 | mipReg; // @[CSR.scala 262:29]
  wire  mip_s_u = _T_2[0]; // @[CSR.scala 262:47]
  wire  mip_s_s = _T_2[1]; // @[CSR.scala 262:47]
  wire  mip_s_h = _T_2[2]; // @[CSR.scala 262:47]
  wire  mip_s_m = _T_2[3]; // @[CSR.scala 262:47]
  wire  mip_t_u = _T_2[4]; // @[CSR.scala 262:47]
  wire  mip_t_s = _T_2[5]; // @[CSR.scala 262:47]
  wire  mip_t_h = _T_2[6]; // @[CSR.scala 262:47]
  wire  mip_t_m = _T_2[7]; // @[CSR.scala 262:47]
  wire  mip_e_u = _T_2[8]; // @[CSR.scala 262:47]
  wire  mip_e_s = _T_2[9]; // @[CSR.scala 262:47]
  wire  mip_e_h = _T_2[10]; // @[CSR.scala 262:47]
  wire  mip_e_m = _T_2[11]; // @[CSR.scala 262:47]
  reg [63:0] misa; // @[CSR.scala 270:21]
  reg [63:0] mstatus; // @[CSR.scala 278:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[CSR.scala 299:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[CSR.scala 299:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[CSR.scala 299:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[CSR.scala 299:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[CSR.scala 299:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[CSR.scala 299:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[CSR.scala 299:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[CSR.scala 299:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[CSR.scala 299:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[CSR.scala 299:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[CSR.scala 299:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[CSR.scala 299:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[CSR.scala 299:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[CSR.scala 299:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[CSR.scala 299:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[CSR.scala 299:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[CSR.scala 299:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[CSR.scala 299:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[CSR.scala 299:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[CSR.scala 299:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[CSR.scala 299:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[CSR.scala 299:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[CSR.scala 299:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[CSR.scala 299:39]
  reg [63:0] medeleg; // @[CSR.scala 306:24]
  reg [63:0] mideleg; // @[CSR.scala 307:24]
  reg [63:0] mscratch; // @[CSR.scala 308:25]
  reg [63:0] pmpcfg0; // @[CSR.scala 310:24]
  reg [63:0] pmpcfg1; // @[CSR.scala 311:24]
  reg [63:0] pmpcfg2; // @[CSR.scala 312:24]
  reg [63:0] pmpcfg3; // @[CSR.scala 313:24]
  reg [63:0] pmpaddr0; // @[CSR.scala 314:25]
  reg [63:0] pmpaddr1; // @[CSR.scala 315:25]
  reg [63:0] pmpaddr2; // @[CSR.scala 316:25]
  reg [63:0] pmpaddr3; // @[CSR.scala 317:25]
  reg [63:0] stvec; // @[CSR.scala 331:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[CSR.scala 333:26]
  reg [63:0] satp; // @[CSR.scala 336:21]
  reg [63:0] sepc; // @[CSR.scala 337:21]
  reg [63:0] scause; // @[CSR.scala 338:23]
  reg [63:0] stval; // @[CSR.scala 339:18]
  reg [63:0] sscratch; // @[CSR.scala 340:25]
  reg [63:0] scounteren; // @[CSR.scala 341:27]
  reg  lr; // @[CSR.scala 354:19]
  reg [63:0] lrAddr; // @[CSR.scala 355:23]
  reg [1:0] priviledgeMode; // @[CSR.scala 368:31]
  reg [63:0] perfCnts_0; // @[CSR.scala 373:47]
  reg [63:0] perfCnts_1; // @[CSR.scala 373:47]
  reg [63:0] perfCnts_2; // @[CSR.scala 373:47]
  wire [5:0] lo_2 = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[CSR.scala 416:27]
  wire [11:0] _T_79 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,lo_2}; // @[CSR.scala 416:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[CSR.scala 456:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[Cat.scala 30:58]
  wire  _T_209 = 12'hf12 == addr; // @[LookupTree.scala 24:34]
  wire  _T_210 = 12'h180 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_247 = _T_210 ? satp : 64'h0; // @[Mux.scala 27:72]
  wire  _T_211 = 12'h3b1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_248 = _T_211 ? pmpaddr1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_284 = _T_247 | _T_248; // @[Mux.scala 27:72]
  wire  _T_212 = 12'h3a2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_249 = _T_212 ? pmpcfg2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_285 = _T_284 | _T_249; // @[Mux.scala 27:72]
  wire  _T_213 = 12'h140 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_250 = _T_213 ? sscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_286 = _T_285 | _T_250; // @[Mux.scala 27:72]
  wire  _T_214 = 12'h302 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_251 = _T_214 ? medeleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_287 = _T_286 | _T_251; // @[Mux.scala 27:72]
  wire  _T_215 = 12'h105 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_252 = _T_215 ? stvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_288 = _T_287 | _T_252; // @[Mux.scala 27:72]
  wire  _T_216 = 12'h141 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_253 = _T_216 ? sepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_289 = _T_288 | _T_253; // @[Mux.scala 27:72]
  wire  _T_217 = 12'h342 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_254 = _T_217 ? mcause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_290 = _T_289 | _T_254; // @[Mux.scala 27:72]
  wire  _T_218 = 12'h306 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_255 = _T_218 ? mcounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_291 = _T_290 | _T_255; // @[Mux.scala 27:72]
  wire  _T_219 = 12'hf11 == addr; // @[LookupTree.scala 24:34]
  wire  _T_220 = 12'h104 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_183 = mie & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_257 = _T_220 ? _T_183 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_293 = _T_291 | _T_257; // @[Mux.scala 27:72]
  wire  _T_221 = 12'h144 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _GEN_79 = {{52'd0}, _T_79}; // @[RegMap.scala 48:84]
  wire [63:0] _T_184 = _GEN_79 & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_258 = _T_221 ? _T_184 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_294 = _T_293 | _T_258; // @[Mux.scala 27:72]
  wire  _T_222 = 12'h100 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_185 = mstatus & 64'h80000003000de122; // @[RegMap.scala 48:84]
  wire [63:0] _T_259 = _T_222 ? _T_185 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_295 = _T_294 | _T_259; // @[Mux.scala 27:72]
  wire  _T_223 = 12'h305 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_260 = _T_223 ? mtvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_296 = _T_295 | _T_260; // @[Mux.scala 27:72]
  wire  _T_224 = 12'h304 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_261 = _T_224 ? mie : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_297 = _T_296 | _T_261; // @[Mux.scala 27:72]
  wire  _T_225 = 12'hb01 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_262 = _T_225 ? perfCnts_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_298 = _T_297 | _T_262; // @[Mux.scala 27:72]
  wire  _T_226 = 12'h3b3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_263 = _T_226 ? pmpaddr3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_299 = _T_298 | _T_263; // @[Mux.scala 27:72]
  wire  _T_227 = 12'h143 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_264 = _T_227 ? stval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_300 = _T_299 | _T_264; // @[Mux.scala 27:72]
  wire  _T_228 = 12'h301 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_265 = _T_228 ? misa : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_301 = _T_300 | _T_265; // @[Mux.scala 27:72]
  wire  _T_229 = 12'h300 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_266 = _T_229 ? mstatus : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_302 = _T_301 | _T_266; // @[Mux.scala 27:72]
  wire  _T_230 = 12'hb00 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_267 = _T_230 ? perfCnts_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_303 = _T_302 | _T_267; // @[Mux.scala 27:72]
  wire  _T_231 = 12'h3b0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_268 = _T_231 ? pmpaddr0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_304 = _T_303 | _T_268; // @[Mux.scala 27:72]
  wire  _T_232 = 12'h344 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_269 = _T_232 ? _GEN_79 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_305 = _T_304 | _T_269; // @[Mux.scala 27:72]
  wire  _T_233 = 12'hb02 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_270 = _T_233 ? perfCnts_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_306 = _T_305 | _T_270; // @[Mux.scala 27:72]
  wire  _T_234 = 12'h3a3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_271 = _T_234 ? pmpcfg3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_307 = _T_306 | _T_271; // @[Mux.scala 27:72]
  wire  _T_235 = 12'h303 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_272 = _T_235 ? mideleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_308 = _T_307 | _T_272; // @[Mux.scala 27:72]
  wire  _T_236 = 12'h3b2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_273 = _T_236 ? pmpaddr2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_309 = _T_308 | _T_273; // @[Mux.scala 27:72]
  wire  _T_237 = 12'hf13 == addr; // @[LookupTree.scala 24:34]
  wire  _T_238 = 12'h3a1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_275 = _T_238 ? pmpcfg1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_311 = _T_309 | _T_275; // @[Mux.scala 27:72]
  wire  _T_239 = 12'h340 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_276 = _T_239 ? mscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_312 = _T_311 | _T_276; // @[Mux.scala 27:72]
  wire  _T_240 = 12'hf14 == addr; // @[LookupTree.scala 24:34]
  wire  _T_241 = 12'h341 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_278 = _T_241 ? mepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_314 = _T_312 | _T_278; // @[Mux.scala 27:72]
  wire  _T_242 = 12'h343 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_279 = _T_242 ? mtval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_315 = _T_314 | _T_279; // @[Mux.scala 27:72]
  wire  _T_243 = 12'h106 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_280 = _T_243 ? scounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_316 = _T_315 | _T_280; // @[Mux.scala 27:72]
  wire  _T_244 = 12'h3a0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_281 = _T_244 ? pmpcfg0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_317 = _T_316 | _T_281; // @[Mux.scala 27:72]
  wire  _T_245 = 12'h142 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_282 = _T_245 ? scause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] rdata = _T_317 | _T_282; // @[Mux.scala 27:72]
  wire [63:0] _T_124 = rdata | io_in_bits_src1; // @[CSR.scala 461:30]
  wire [63:0] _T_125 = ~io_in_bits_src1; // @[CSR.scala 462:32]
  wire [63:0] _T_126 = rdata & _T_125; // @[CSR.scala 462:30]
  wire [63:0] _T_127 = rdata | csri; // @[CSR.scala 464:30]
  wire [63:0] _T_128 = ~csri; // @[CSR.scala 465:32]
  wire [63:0] _T_129 = rdata & _T_128; // @[CSR.scala 465:30]
  wire  _T_130 = 7'h1 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_131 = 7'h2 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_132 = 7'h3 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_133 = 7'h5 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_134 = 7'h6 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_135 = 7'h7 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_136 = _T_130 ? io_in_bits_src1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_137 = _T_131 ? _T_124 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_138 = _T_132 ? _T_126 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_139 = _T_133 ? csri : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_140 = _T_134 ? _T_127 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_141 = _T_135 ? _T_129 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_142 = _T_136 | _T_137; // @[Mux.scala 27:72]
  wire [63:0] _T_143 = _T_142 | _T_138; // @[Mux.scala 27:72]
  wire [63:0] _T_144 = _T_143 | _T_139; // @[Mux.scala 27:72]
  wire [63:0] _T_145 = _T_144 | _T_140; // @[Mux.scala 27:72]
  wire [63:0] wdata = _T_145 | _T_141; // @[Mux.scala 27:72]
  wire  satpLegalMode = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[CSR.scala 469:69]
  wire  wen = io_in_valid & io_in_bits_func != 7'h0 & (addr != 12'h180 | satpLegalMode); // @[CSR.scala 472:47]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[CSR.scala 473:39]
  wire  justRead = (io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6) & io_in_bits_src1 == 64'h0; // @[CSR.scala 474:70]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~justRead; // @[CSR.scala 475:58]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite; // @[CSR.scala 476:39]
  wire  _T_171 = wen & ~isIllegalAccess; // @[CSR.scala 478:51]
  wire  _T_319 = addr == 12'h180; // @[RegMap.scala 50:65]
  wire  _T_343 = addr == 12'h302; // @[RegMap.scala 50:65]
  wire [63:0] _T_345 = wdata & 64'hbbff; // @[BitUtils.scala 32:13]
  wire [63:0] _T_347 = medeleg & 64'h4400; // @[BitUtils.scala 32:36]
  wire [63:0] _T_348 = _T_345 | _T_347; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_8 = _T_171 & addr == 12'h141 ? wdata : sepc; // @[CSR.scala 337:21 RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_9 = _T_171 & addr == 12'h342 ? wdata : mcause; // @[CSR.scala 254:23 RegMap.scala 50:{72,76}]
  wire [63:0] _T_375 = wdata & sieMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_376 = ~sieMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_377 = mie & _T_376; // @[BitUtils.scala 32:36]
  wire [63:0] _T_378 = _T_375 | _T_377; // @[BitUtils.scala 32:25]
  wire [63:0] _T_381 = wdata & 64'hc6122; // @[BitUtils.scala 32:13]
  wire [63:0] _T_383 = mstatus & 64'h39edd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_384 = _T_381 | _T_383; // @[BitUtils.scala 32:25]
  wire  _T_409 = _T_384[14:13] == 2'h3; // @[CSR.scala 302:40]
  wire [63:0] _T_411 = {_T_409,_T_384[62:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_12 = _T_171 & addr == 12'h100 ? _T_411 : mstatus; // @[CSR.scala 278:24 RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_17 = _T_171 & addr == 12'h143 ? wdata : stval; // @[CSR.scala 339:18 RegMap.scala 50:{72,76}]
  wire  _T_478 = wdata[14:13] == 2'h3; // @[CSR.scala 302:40]
  wire [63:0] _T_480 = {_T_478,wdata[62:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_19 = _T_171 & addr == 12'h300 ? _T_480 : _GEN_12; // @[RegMap.scala 50:{72,76}]
  wire [63:0] _T_507 = wdata & 64'h222; // @[BitUtils.scala 32:13]
  wire [63:0] _T_509 = mideleg & 64'h1dd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_510 = _T_507 | _T_509; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_28 = _T_171 & addr == 12'h341 ? wdata : mepc; // @[CSR.scala 256:17 RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_29 = _T_171 & addr == 12'h343 ? wdata : mtval; // @[CSR.scala 255:22 RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_32 = _T_171 & addr == 12'h142 ? wdata : scause; // @[CSR.scala 338:23 RegMap.scala 50:{72,76}]
  wire  _T_560 = _T_209 ? 1'h0 : 1'h1; // @[Mux.scala 80:57]
  wire  _T_562 = _T_210 ? 1'h0 : _T_560; // @[Mux.scala 80:57]
  wire  _T_564 = _T_211 ? 1'h0 : _T_562; // @[Mux.scala 80:57]
  wire  _T_566 = _T_212 ? 1'h0 : _T_564; // @[Mux.scala 80:57]
  wire  _T_568 = _T_213 ? 1'h0 : _T_566; // @[Mux.scala 80:57]
  wire  _T_570 = _T_214 ? 1'h0 : _T_568; // @[Mux.scala 80:57]
  wire  _T_572 = _T_215 ? 1'h0 : _T_570; // @[Mux.scala 80:57]
  wire  _T_574 = _T_216 ? 1'h0 : _T_572; // @[Mux.scala 80:57]
  wire  _T_576 = _T_217 ? 1'h0 : _T_574; // @[Mux.scala 80:57]
  wire  _T_578 = _T_218 ? 1'h0 : _T_576; // @[Mux.scala 80:57]
  wire  _T_580 = _T_219 ? 1'h0 : _T_578; // @[Mux.scala 80:57]
  wire  _T_582 = _T_220 ? 1'h0 : _T_580; // @[Mux.scala 80:57]
  wire  _T_584 = _T_221 ? 1'h0 : _T_582; // @[Mux.scala 80:57]
  wire  _T_586 = _T_222 ? 1'h0 : _T_584; // @[Mux.scala 80:57]
  wire  _T_588 = _T_223 ? 1'h0 : _T_586; // @[Mux.scala 80:57]
  wire  _T_590 = _T_224 ? 1'h0 : _T_588; // @[Mux.scala 80:57]
  wire  _T_592 = _T_225 ? 1'h0 : _T_590; // @[Mux.scala 80:57]
  wire  _T_594 = _T_226 ? 1'h0 : _T_592; // @[Mux.scala 80:57]
  wire  _T_596 = _T_227 ? 1'h0 : _T_594; // @[Mux.scala 80:57]
  wire  _T_598 = _T_228 ? 1'h0 : _T_596; // @[Mux.scala 80:57]
  wire  _T_600 = _T_229 ? 1'h0 : _T_598; // @[Mux.scala 80:57]
  wire  _T_602 = _T_230 ? 1'h0 : _T_600; // @[Mux.scala 80:57]
  wire  _T_604 = _T_231 ? 1'h0 : _T_602; // @[Mux.scala 80:57]
  wire  _T_606 = _T_232 ? 1'h0 : _T_604; // @[Mux.scala 80:57]
  wire  _T_608 = _T_233 ? 1'h0 : _T_606; // @[Mux.scala 80:57]
  wire  _T_610 = _T_234 ? 1'h0 : _T_608; // @[Mux.scala 80:57]
  wire  _T_612 = _T_235 ? 1'h0 : _T_610; // @[Mux.scala 80:57]
  wire  _T_614 = _T_236 ? 1'h0 : _T_612; // @[Mux.scala 80:57]
  wire  _T_616 = _T_237 ? 1'h0 : _T_614; // @[Mux.scala 80:57]
  wire  _T_618 = _T_238 ? 1'h0 : _T_616; // @[Mux.scala 80:57]
  wire  _T_620 = _T_239 ? 1'h0 : _T_618; // @[Mux.scala 80:57]
  wire  _T_622 = _T_240 ? 1'h0 : _T_620; // @[Mux.scala 80:57]
  wire  _T_624 = _T_241 ? 1'h0 : _T_622; // @[Mux.scala 80:57]
  wire  _T_626 = _T_242 ? 1'h0 : _T_624; // @[Mux.scala 80:57]
  wire  _T_628 = _T_243 ? 1'h0 : _T_626; // @[Mux.scala 80:57]
  wire  _T_630 = _T_244 ? 1'h0 : _T_628; // @[Mux.scala 80:57]
  wire  isIllegalAddr = _T_245 ? 1'h0 : _T_630; // @[Mux.scala 80:57]
  wire  resetSatp = _T_319 & wen; // @[CSR.scala 480:35]
  wire [63:0] _T_646 = wdata & 64'h77f; // @[BitUtils.scala 32:13]
  wire [63:0] _T_648 = mipReg & 64'h80; // @[BitUtils.scala 32:36]
  wire [63:0] _T_649 = _T_646 | _T_648; // @[BitUtils.scala 32:25]
  wire [63:0] _T_654 = mipReg & _T_376; // @[BitUtils.scala 32:36]
  wire [63:0] _T_655 = _T_375 | _T_654; // @[BitUtils.scala 32:25]
  wire  _T_657 = io_in_bits_func == 7'h0; // @[CSR.scala 493:46]
  wire  isEbreak = addr == 12'h1 & io_in_bits_func == 7'h0; // @[CSR.scala 493:38]
  wire  isEcall = addr == 12'h0 & _T_657; // @[CSR.scala 494:36]
  wire  isMret = _T_343 & _T_657; // @[CSR.scala 495:36]
  wire  isSret = addr == 12'h102 & _T_657; // @[CSR.scala 496:36]
  wire  isUret = addr == 12'h2 & _T_657; // @[CSR.scala 497:36]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_in_valid; // @[CSR.scala 554:63]
  wire  _T_699 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF; // @[CSR.scala 563:46]
  wire [38:0] _T_701 = io_cfIn_pc + 39'h2; // @[CSR.scala 564:88]
  wire [24:0] _T_705 = _T_701[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_706 = {_T_705,_T_701}; // @[Cat.scala 30:58]
  wire [24:0] _T_710 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_711 = {_T_710,io_cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_712 = io_cfIn_crossPageIPFFix ? _T_706 : _T_711; // @[CSR.scala 564:42]
  wire [24:0] _T_715 = io_dmemMMU_addr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_716 = {_T_715,io_dmemMMU_addr}; // @[Cat.scala 30:58]
  wire [63:0] _T_717 = hasInstrPageFault ? _T_712 : _T_716; // @[CSR.scala 564:19]
  wire  _T_718 = priviledgeMode == 2'h3; // @[CSR.scala 565:25]
  wire [63:0] _GEN_35 = priviledgeMode == 2'h3 ? _T_717 : _GEN_29; // @[CSR.scala 565:35 566:13]
  wire [63:0] _GEN_36 = priviledgeMode == 2'h3 ? _GEN_17 : _T_717; // @[CSR.scala 565:35 568:13]
  wire [63:0] _GEN_37 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF ? _GEN_35 : _GEN_29; // @[CSR.scala 563:67]
  wire [63:0] _GEN_38 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF ? _GEN_36 : _GEN_17; // @[CSR.scala 563:67]
  wire  _T_732 = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[CSR.scala 573:30]
  wire [38:0] dmemAddrMisalignedAddr = LSUADDR[38:0]; // @[CSR.scala 542:36 560:28]
  wire [24:0] _T_735 = dmemAddrMisalignedAddr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_736 = {_T_735,dmemAddrMisalignedAddr}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_39 = _T_732 ? _T_736 : _GEN_37; // @[CSR.scala 574:3 575:11]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[CSR.scala 597:31]
  wire [11:0] _T_751 = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,lo_2}; // @[CSR.scala 599:41]
  wire [63:0] _GEN_80 = {{52'd0}, _T_751}; // @[CSR.scala 599:26]
  wire [63:0] ideleg = mideleg & _GEN_80; // @[CSR.scala 599:26]
  wire  _T_816 = priviledgeMode == 2'h1; // @[CSR.scala 600:72]
  wire  _T_822 = priviledgeMode < 2'h3; // @[CSR.scala 601:106]
  wire  _T_823 = _T_718 & mstatusStruct_ie_m | priviledgeMode < 2'h3; // @[CSR.scala 601:87]
  wire  intrVecEnable_0 = ideleg[0] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_1 = ideleg[1] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_2 = ideleg[2] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_3 = ideleg[3] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_4 = ideleg[4] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_5 = ideleg[5] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_6 = ideleg[6] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_7 = ideleg[7] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_8 = ideleg[8] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_9 = ideleg[9] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_10 = ideleg[10] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire  intrVecEnable_11 = ideleg[11] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_823; // @[CSR.scala 600:51]
  wire [11:0] _T_926 = mie[11:0] & _T_751; // @[CSR.scala 605:27]
  wire [5:0] lo_6 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,intrVecEnable_0}; // @[CSR.scala 605:65]
  wire [11:0] _T_927 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,lo_6}; // @[CSR.scala 605:65]
  wire [11:0] intrVec = _T_926 & _T_927; // @[CSR.scala 605:49]
  wire [2:0] _T_928 = io_cfIn_intrVec_4 ? 3'h4 : 3'h0; // @[CSR.scala 609:69]
  wire [3:0] _T_929 = io_cfIn_intrVec_8 ? 4'h8 : {{1'd0}, _T_928}; // @[CSR.scala 609:69]
  wire [3:0] _T_930 = io_cfIn_intrVec_0 ? 4'h0 : _T_929; // @[CSR.scala 609:69]
  wire [3:0] _T_931 = io_cfIn_intrVec_5 ? 4'h5 : _T_930; // @[CSR.scala 609:69]
  wire [3:0] _T_932 = io_cfIn_intrVec_9 ? 4'h9 : _T_931; // @[CSR.scala 609:69]
  wire [3:0] _T_933 = io_cfIn_intrVec_1 ? 4'h1 : _T_932; // @[CSR.scala 609:69]
  wire [3:0] _T_934 = io_cfIn_intrVec_7 ? 4'h7 : _T_933; // @[CSR.scala 609:69]
  wire [3:0] _T_935 = io_cfIn_intrVec_11 ? 4'hb : _T_934; // @[CSR.scala 609:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _T_935; // @[CSR.scala 609:69]
  wire [5:0] lo_7 = {io_cfIn_intrVec_5,io_cfIn_intrVec_4,io_cfIn_intrVec_3,io_cfIn_intrVec_2,io_cfIn_intrVec_1,
    io_cfIn_intrVec_0}; // @[CSR.scala 611:35]
  wire [11:0] _T_936 = {io_cfIn_intrVec_11,io_cfIn_intrVec_10,io_cfIn_intrVec_9,io_cfIn_intrVec_8,io_cfIn_intrVec_7,
    io_cfIn_intrVec_6,lo_7}; // @[CSR.scala 611:35]
  wire  raiseIntr = |_T_936; // @[CSR.scala 611:42]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[CSR.scala 618:46]
  wire  csrExceptionVec_11 = _T_718 & io_in_valid & isEcall; // @[CSR.scala 619:70]
  wire  csrExceptionVec_9 = _T_816 & io_in_valid & isEcall; // @[CSR.scala 620:70]
  wire  csrExceptionVec_8 = priviledgeMode == 2'h0 & io_in_valid & isEcall; // @[CSR.scala 621:70]
  wire  csrExceptionVec_2 = (isIllegalAddr | isIllegalAccess) & wen; // @[CSR.scala 622:71]
  wire [7:0] lo_8 = {4'h0,csrExceptionVec_3,csrExceptionVec_2,2'h0}; // @[CSR.scala 626:49]
  wire [15:0] _T_951 = {io_dmemMMU_storePF,1'h0,io_dmemMMU_loadPF,1'h0,csrExceptionVec_11,1'h0,csrExceptionVec_9,
    csrExceptionVec_8,lo_8}; // @[CSR.scala 626:49]
  wire [7:0] lo_9 = {1'h0,io_cfIn_exceptionVec_6,1'h0,io_cfIn_exceptionVec_4,1'h0,io_cfIn_exceptionVec_2,
    io_cfIn_exceptionVec_1,1'h0}; // @[CSR.scala 626:76]
  wire [15:0] _T_952 = {2'h0,1'h0,io_cfIn_exceptionVec_12,4'h0,lo_9}; // @[CSR.scala 626:76]
  wire [15:0] raiseExceptionVec = _T_951 | _T_952; // @[CSR.scala 626:52]
  wire  raiseException = |raiseExceptionVec; // @[CSR.scala 627:42]
  wire [2:0] _T_954 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[CSR.scala 628:74]
  wire [2:0] _T_956 = raiseExceptionVec[7] ? 3'h7 : _T_954; // @[CSR.scala 628:74]
  wire [3:0] _T_958 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _T_956}; // @[CSR.scala 628:74]
  wire [3:0] _T_960 = raiseExceptionVec[15] ? 4'hf : _T_958; // @[CSR.scala 628:74]
  wire [3:0] _T_962 = raiseExceptionVec[4] ? 4'h4 : _T_960; // @[CSR.scala 628:74]
  wire [3:0] _T_964 = raiseExceptionVec[6] ? 4'h6 : _T_962; // @[CSR.scala 628:74]
  wire [3:0] _T_966 = raiseExceptionVec[8] ? 4'h8 : _T_964; // @[CSR.scala 628:74]
  wire [3:0] _T_968 = raiseExceptionVec[9] ? 4'h9 : _T_966; // @[CSR.scala 628:74]
  wire [3:0] _T_970 = raiseExceptionVec[11] ? 4'hb : _T_968; // @[CSR.scala 628:74]
  wire [3:0] _T_972 = raiseExceptionVec[0] ? 4'h0 : _T_970; // @[CSR.scala 628:74]
  wire [3:0] _T_974 = raiseExceptionVec[2] ? 4'h2 : _T_972; // @[CSR.scala 628:74]
  wire [3:0] _T_976 = raiseExceptionVec[1] ? 4'h1 : _T_974; // @[CSR.scala 628:74]
  wire [3:0] _T_978 = raiseExceptionVec[12] ? 4'hc : _T_976; // @[CSR.scala 628:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _T_978; // @[CSR.scala 628:74]
  wire [63:0] _T_980 = {raiseIntr, 63'h0}; // @[CSR.scala 631:28]
  wire [3:0] _T_981 = raiseIntr ? intrNO : exceptionNO; // @[CSR.scala 631:46]
  wire [63:0] _GEN_81 = {{60'd0}, _T_981}; // @[CSR.scala 631:41]
  wire [63:0] causeNO = _T_980 | _GEN_81; // @[CSR.scala 631:41]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid; // @[CSR.scala 634:58]
  wire [38:0] _T_989 = io_cfIn_pc + 39'h4; // @[CSR.scala 639:51]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[CSR.scala 649:18]
  wire [63:0] _T_1033 = deleg >> causeNO[3:0]; // @[CSR.scala 651:22]
  wire  delegS = _T_1033[0] & _T_822; // @[CSR.scala 651:38]
  wire [63:0] _T_1043 = delegS ? stvec : mtvec; // @[CSR.scala 655:20]
  wire [38:0] trapTarget = _T_1043[38:0]; // @[CSR.scala 655:42]
  wire [38:0] _GEN_47 = io_in_valid & isSret ? sepc[38:0] : mepc[38:0]; // @[CSR.scala 673:26 683:15]
  wire [38:0] retTarget = io_in_valid & isUret ? 39'h0 : _GEN_47; // @[CSR.scala 686:26 694:15]
  wire [38:0] _T_990 = raiseExceptionIntr ? trapTarget : retTarget; // @[CSR.scala 639:61]
  wire  tvalWen = ~(_T_699 | io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6) | raiseIntr; // @[CSR.scala 652:130]
  wire [5:0] lo_lo_13 = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,
    mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[CSR.scala 668:27]
  wire [14:0] lo_13 = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,lo_lo_13}; // @[CSR.scala 668:27]
  wire [6:0] hi_lo_13 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusStruct_mprv,
    mstatusStruct_xs}; // @[CSR.scala 668:27]
  wire [63:0] _T_1094 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_13,lo_13}; // @[CSR.scala 668:27]
  wire [1:0] _GEN_40 = io_in_valid & isMret ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 660:26 665:20 368:31]
  wire [63:0] _GEN_41 = io_in_valid & isMret ? _T_1094 : _GEN_19; // @[CSR.scala 660:26 668:13]
  wire [1:0] _T_1145 = {1'h0,mstatusStruct_spp}; // @[Cat.scala 30:58]
  wire [5:0] lo_lo_14 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,
    mstatusStruct_ie_u}; // @[CSR.scala 681:27]
  wire [14:0] lo_14 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,mstatusStruct_pie_h
    ,lo_lo_14}; // @[CSR.scala 681:27]
  wire [63:0] _T_1146 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_13,lo_14}; // @[CSR.scala 681:27]
  wire [5:0] lo_lo_15 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,
    mstatusStruct_pie_u}; // @[CSR.scala 693:27]
  wire [14:0] lo_15 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m,
    mstatusStruct_pie_h,lo_lo_15}; // @[CSR.scala 693:27]
  wire [63:0] _T_1197 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_13,lo_15}; // @[CSR.scala 693:27]
  wire [1:0] _GEN_55 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[CSR.scala 701:19 704:22]
  wire  _GEN_56 = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[CSR.scala 701:19 705:24]
  wire  _GEN_57 = delegS ? 1'h0 : mstatusStruct_ie_s; // @[CSR.scala 701:19 706:23]
  wire [1:0] _GEN_62 = delegS ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 701:19 714:22]
  wire  _GEN_63 = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[CSR.scala 701:19 715:24]
  wire  _GEN_64 = delegS & mstatusStruct_ie_m; // @[CSR.scala 701:19 716:23]
  wire [5:0] lo_lo_16 = {_GEN_56,mstatusStruct_pie_u,_GEN_64,mstatusStruct_ie_h,_GEN_57,mstatusStruct_ie_u}; // @[CSR.scala 728:27]
  wire [14:0] lo_16 = {mstatusStruct_fs,_GEN_62,mstatusStruct_hpp,_GEN_55[0],_GEN_63,mstatusStruct_pie_h,lo_lo_16}; // @[CSR.scala 728:27]
  wire [63:0] _T_1255 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_13,lo_16}; // @[CSR.scala 728:27]
  wire [63:0] _T_1257 = perfCnts_0 + 64'h1; // @[CSR.scala 837:71]
  wire  _WIRE_49 = 1'h1;
  wire [63:0] _T_1261 = perfCnts_2 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_1263 = perfCnts_2 + 64'h2; // @[CSR.scala 845:86]
  assign io_out_valid = io_in_valid; // @[CSR.scala 732:16]
  assign io_out_bits = _T_317 | _T_282; // @[Mux.scala 27:72]
  assign io_redirect_target = resetSatp ? _T_989 : _T_990; // @[CSR.scala 639:28]
  assign io_redirect_valid = io_in_valid & _T_657 | raiseExceptionIntr | resetSatp; // @[CSR.scala 637:80]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[CSR.scala 528:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 529:35]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[CSR.scala 299:39]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[CSR.scala 299:39]
  assign io_wenFix = |raiseExceptionVec; // @[CSR.scala 627:42]
  assign perfCnts_2_0 = perfCnts_2;
  assign satp_0 = satp;
  assign intrVec_0 = intrVec;
  assign lrAddr_0 = lrAddr;
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 252:22]
      mtvec <= 64'h0; // @[CSR.scala 252:22]
    end else if (_T_171 & addr == 12'h305) begin // @[RegMap.scala 50:72]
      mtvec <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 253:27]
      mcounteren <= 64'h0; // @[CSR.scala 253:27]
    end else if (_T_171 & addr == 12'h306) begin // @[RegMap.scala 50:72]
      mcounteren <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 254:23]
      mcause <= 64'h0; // @[CSR.scala 254:23]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      if (delegS) begin // @[CSR.scala 701:19]
        mcause <= _GEN_9;
      end else begin
        mcause <= causeNO; // @[CSR.scala 712:14]
      end
    end else begin
      mcause <= _GEN_9;
    end
    if (reset) begin // @[CSR.scala 255:22]
      mtval <= 64'h0; // @[CSR.scala 255:22]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      if (delegS) begin // @[CSR.scala 701:19]
        mtval <= _GEN_39;
      end else if (tvalWen) begin // @[CSR.scala 718:20]
        mtval <= 64'h0; // @[CSR.scala 718:27]
      end else begin
        mtval <= _GEN_39;
      end
    end else begin
      mtval <= _GEN_39;
    end
    if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      if (delegS) begin // @[CSR.scala 701:19]
        mepc <= _GEN_28;
      end else begin
        mepc <= _T_711; // @[CSR.scala 713:12]
      end
    end else begin
      mepc <= _GEN_28;
    end
    if (reset) begin // @[CSR.scala 258:20]
      mie <= 64'h0; // @[CSR.scala 258:20]
    end else if (_T_171 & addr == 12'h304) begin // @[RegMap.scala 50:72]
      mie <= wdata; // @[RegMap.scala 50:76]
    end else if (_T_171 & addr == 12'h104) begin // @[RegMap.scala 50:72]
      mie <= _T_378; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 260:24]
      mipReg <= 64'h0; // @[CSR.scala 260:24]
    end else if (_T_171 & addr == 12'h144) begin // @[RegMap.scala 50:72]
      mipReg <= _T_655; // @[RegMap.scala 50:76]
    end else if (_T_171 & addr == 12'h344) begin // @[RegMap.scala 50:72]
      mipReg <= _T_649; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 270:21]
      misa <= 64'h8000000000141105; // @[CSR.scala 270:21]
    end else if (_T_171 & addr == 12'h301) begin // @[RegMap.scala 50:72]
      misa <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 278:24]
      mstatus <= 64'h1800; // @[CSR.scala 278:24]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      mstatus <= _T_1255; // @[CSR.scala 728:13]
    end else if (io_in_valid & isUret) begin // @[CSR.scala 686:26]
      mstatus <= _T_1197; // @[CSR.scala 693:13]
    end else if (io_in_valid & isSret) begin // @[CSR.scala 673:26]
      mstatus <= _T_1146; // @[CSR.scala 681:13]
    end else begin
      mstatus <= _GEN_41;
    end
    if (reset) begin // @[CSR.scala 306:24]
      medeleg <= 64'h0; // @[CSR.scala 306:24]
    end else if (_T_171 & addr == 12'h302) begin // @[RegMap.scala 50:72]
      medeleg <= _T_348; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 307:24]
      mideleg <= 64'h0; // @[CSR.scala 307:24]
    end else if (_T_171 & addr == 12'h303) begin // @[RegMap.scala 50:72]
      mideleg <= _T_510; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 308:25]
      mscratch <= 64'h0; // @[CSR.scala 308:25]
    end else if (_T_171 & addr == 12'h340) begin // @[RegMap.scala 50:72]
      mscratch <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 310:24]
      pmpcfg0 <= 64'h0; // @[CSR.scala 310:24]
    end else if (_T_171 & addr == 12'h3a0) begin // @[RegMap.scala 50:72]
      pmpcfg0 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 311:24]
      pmpcfg1 <= 64'h0; // @[CSR.scala 311:24]
    end else if (_T_171 & addr == 12'h3a1) begin // @[RegMap.scala 50:72]
      pmpcfg1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 312:24]
      pmpcfg2 <= 64'h0; // @[CSR.scala 312:24]
    end else if (_T_171 & addr == 12'h3a2) begin // @[RegMap.scala 50:72]
      pmpcfg2 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 313:24]
      pmpcfg3 <= 64'h0; // @[CSR.scala 313:24]
    end else if (_T_171 & addr == 12'h3a3) begin // @[RegMap.scala 50:72]
      pmpcfg3 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 314:25]
      pmpaddr0 <= 64'h0; // @[CSR.scala 314:25]
    end else if (_T_171 & addr == 12'h3b0) begin // @[RegMap.scala 50:72]
      pmpaddr0 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 315:25]
      pmpaddr1 <= 64'h0; // @[CSR.scala 315:25]
    end else if (_T_171 & addr == 12'h3b1) begin // @[RegMap.scala 50:72]
      pmpaddr1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 316:25]
      pmpaddr2 <= 64'h0; // @[CSR.scala 316:25]
    end else if (_T_171 & addr == 12'h3b2) begin // @[RegMap.scala 50:72]
      pmpaddr2 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 317:25]
      pmpaddr3 <= 64'h0; // @[CSR.scala 317:25]
    end else if (_T_171 & addr == 12'h3b3) begin // @[RegMap.scala 50:72]
      pmpaddr3 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 331:22]
      stvec <= 64'h0; // @[CSR.scala 331:22]
    end else if (_T_171 & addr == 12'h105) begin // @[RegMap.scala 50:72]
      stvec <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 336:21]
      satp <= 64'h0; // @[CSR.scala 336:21]
    end else if (_T_171 & addr == 12'h180) begin // @[RegMap.scala 50:72]
      satp <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 337:21]
      sepc <= 64'h0; // @[CSR.scala 337:21]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      if (delegS) begin // @[CSR.scala 701:19]
        sepc <= _T_711; // @[CSR.scala 703:12]
      end else begin
        sepc <= _GEN_8;
      end
    end else begin
      sepc <= _GEN_8;
    end
    if (reset) begin // @[CSR.scala 338:23]
      scause <= 64'h0; // @[CSR.scala 338:23]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      if (delegS) begin // @[CSR.scala 701:19]
        scause <= causeNO; // @[CSR.scala 702:14]
      end else begin
        scause <= _GEN_32;
      end
    end else begin
      scause <= _GEN_32;
    end
    if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      if (delegS) begin // @[CSR.scala 701:19]
        if (tvalWen) begin // @[CSR.scala 708:20]
          stval <= 64'h0; // @[CSR.scala 708:27]
        end else begin
          stval <= _GEN_38;
        end
      end else begin
        stval <= _GEN_38;
      end
    end else begin
      stval <= _GEN_38;
    end
    if (reset) begin // @[CSR.scala 340:25]
      sscratch <= 64'h0; // @[CSR.scala 340:25]
    end else if (_T_171 & addr == 12'h140) begin // @[RegMap.scala 50:72]
      sscratch <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 341:27]
      scounteren <= 64'h0; // @[CSR.scala 341:27]
    end else if (_T_171 & addr == 12'h106) begin // @[RegMap.scala 50:72]
      scounteren <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 354:19]
      lr <= 1'h0; // @[CSR.scala 354:19]
    end else if (io_in_valid & isSret) begin // @[CSR.scala 673:26]
      lr <= 1'h0; // @[CSR.scala 682:8]
    end else if (io_in_valid & isMret) begin // @[CSR.scala 660:26]
      lr <= 1'h0; // @[CSR.scala 669:8]
    end else if (set_lr) begin // @[CSR.scala 362:14]
      lr <= set_lr_val; // @[CSR.scala 363:8]
    end
    if (reset) begin // @[CSR.scala 355:23]
      lrAddr <= 64'h0; // @[CSR.scala 355:23]
    end else if (set_lr) begin // @[CSR.scala 362:14]
      lrAddr <= set_lr_addr; // @[CSR.scala 364:12]
    end
    if (reset) begin // @[CSR.scala 368:31]
      priviledgeMode <= 2'h3; // @[CSR.scala 368:31]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 697:29]
      if (delegS) begin // @[CSR.scala 701:19]
        priviledgeMode <= 2'h1; // @[CSR.scala 707:22]
      end else begin
        priviledgeMode <= 2'h3; // @[CSR.scala 717:22]
      end
    end else if (io_in_valid & isUret) begin // @[CSR.scala 686:26]
      priviledgeMode <= 2'h0; // @[CSR.scala 691:20]
    end else if (io_in_valid & isSret) begin // @[CSR.scala 673:26]
      priviledgeMode <= _T_1145; // @[CSR.scala 678:20]
    end else begin
      priviledgeMode <= _GEN_40;
    end
    if (reset) begin // @[CSR.scala 373:47]
      perfCnts_0 <= 64'h0; // @[CSR.scala 373:47]
    end else begin
      perfCnts_0 <= _T_1257;
    end
    if (reset) begin // @[CSR.scala 373:47]
      perfCnts_1 <= 64'h0; // @[CSR.scala 373:47]
    end else if (_T_171 & addr == 12'hb01) begin // @[RegMap.scala 50:72]
      perfCnts_1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 373:47]
      perfCnts_2 <= 64'h0; // @[CSR.scala 373:47]
    end else if (perfCntCondMultiCommit) begin // @[CSR.scala 845:35]
      perfCnts_2 <= _T_1263; // @[CSR.scala 845:60]
    end else if (perfCntCondMinstret) begin // @[CSR.scala 837:62]
      perfCnts_2 <= _T_1261; // @[CSR.scala 837:66]
    end else if (_T_171 & addr == 12'hb02) begin // @[RegMap.scala 50:72]
      perfCnts_2 <= wdata; // @[RegMap.scala 50:76]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtval = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mipReg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  misa = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  pmpcfg0 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pmpcfg1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  pmpcfg2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  pmpcfg3 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  pmpaddr0 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  pmpaddr1 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  pmpaddr2 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  pmpaddr3 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  stvec = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  satp = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  sepc = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  scause = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  stval = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  sscratch = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  scounteren = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  lr = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  lrAddr = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  priviledgeMode = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  perfCnts_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  perfCnts_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  perfCnts_2 = _RAND_32[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MOU(
  input         io_in_valid,
  input  [6:0]  io_in_bits_func,
  input  [38:0] io_cfIn_pc,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  output        flushICache_0,
  output        flushTLB_0
);
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1; // @[MOU.scala 52:27]
  wire  flushTLB = io_in_valid & io_in_bits_func == 7'h2; // @[MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[MOU.scala 49:36]
  assign io_redirect_valid = io_in_valid; // @[MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io__in_ready,
  input         io__in_valid,
  input  [63:0] io__in_bits_cf_instr,
  input  [38:0] io__in_bits_cf_pc,
  input  [38:0] io__in_bits_cf_pnpc,
  input         io__in_bits_cf_exceptionVec_1,
  input         io__in_bits_cf_exceptionVec_2,
  input         io__in_bits_cf_exceptionVec_12,
  input         io__in_bits_cf_intrVec_0,
  input         io__in_bits_cf_intrVec_1,
  input         io__in_bits_cf_intrVec_2,
  input         io__in_bits_cf_intrVec_3,
  input         io__in_bits_cf_intrVec_4,
  input         io__in_bits_cf_intrVec_5,
  input         io__in_bits_cf_intrVec_6,
  input         io__in_bits_cf_intrVec_7,
  input         io__in_bits_cf_intrVec_8,
  input         io__in_bits_cf_intrVec_9,
  input         io__in_bits_cf_intrVec_10,
  input         io__in_bits_cf_intrVec_11,
  input  [3:0]  io__in_bits_cf_brIdx,
  input         io__in_bits_cf_crossPageIPFFix,
  input  [63:0] io__in_bits_cf_runahead_checkpoint_id,
  input  [2:0]  io__in_bits_ctrl_fuType,
  input  [6:0]  io__in_bits_ctrl_fuOpType,
  input         io__in_bits_ctrl_rfWen,
  input  [4:0]  io__in_bits_ctrl_rfDest,
  input  [2:0]  io__in_bits_ctrl_vtag,
  input  [4:0]  io__in_bits_ctrl_vec_addr,
  input  [3:0]  io__in_bits_ctrl_length_k,
  input  [1:0]  io__in_bits_ctrl_algorithm,
  input  [63:0] io__in_bits_data_src1,
  input  [63:0] io__in_bits_data_src2,
  input  [63:0] io__in_bits_data_imm,
  input         io__out_ready,
  output        io__out_valid,
  output [38:0] io__out_bits_decode_cf_pc,
  output [38:0] io__out_bits_decode_cf_redirect_target,
  output        io__out_bits_decode_cf_redirect_valid,
  output [63:0] io__out_bits_decode_cf_runahead_checkpoint_id,
  output [2:0]  io__out_bits_decode_ctrl_fuType,
  output        io__out_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_bits_decode_ctrl_rfDest,
  output [63:0] io__out_bits_commits_0,
  output [63:0] io__out_bits_commits_1,
  output [63:0] io__out_bits_commits_2,
  output [63:0] io__out_bits_commits_3,
  output [63:0] io__out_bits_commits_5,
  input         io__flush,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__forward_valid,
  output        io__forward_wb_rfWen,
  output [4:0]  io__forward_wb_rfDest,
  output [63:0] io__forward_wb_rfData,
  output [2:0]  io__forward_fuType,
  output [1:0]  io__memMMU_imem_priviledgeMode,
  output [1:0]  io__memMMU_dmem_priviledgeMode,
  output        io__memMMU_dmem_status_sum,
  output        io__memMMU_dmem_status_mxr,
  input         io__memMMU_dmem_loadPF,
  input         io__memMMU_dmem_storePF,
  input  [38:0] io__memMMU_dmem_addr,
  input         _T_28_0,
  output        flushICache,
  output [63:0] perfCnts_2,
  output [63:0] satp,
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output        REG_0_actualTaken,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC,
  input         io_in_valid,
  input         io_extra_mtip,
  output        amoReq,
  input         io_extra_meip_0,
  input         vmEnable,
  output [11:0] intrVec,
  input         _T_27_0,
  input         io_extra_msip,
  output        flushTLB,
  input         falseWire
);
  wire  alu_clock; // @[EXU.scala 48:19]
  wire  alu_reset; // @[EXU.scala 48:19]
  wire  alu_io_in_valid; // @[EXU.scala 48:19]
  wire [63:0] alu_io_in_bits_src1; // @[EXU.scala 48:19]
  wire [63:0] alu_io_in_bits_src2; // @[EXU.scala 48:19]
  wire [6:0] alu_io_in_bits_func; // @[EXU.scala 48:19]
  wire  alu_io_out_ready; // @[EXU.scala 48:19]
  wire  alu_io_out_valid; // @[EXU.scala 48:19]
  wire [63:0] alu_io_out_bits; // @[EXU.scala 48:19]
  wire [63:0] alu_io_cfIn_instr; // @[EXU.scala 48:19]
  wire [38:0] alu_io_cfIn_pc; // @[EXU.scala 48:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[EXU.scala 48:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[EXU.scala 48:19]
  wire [38:0] alu_io_redirect_target; // @[EXU.scala 48:19]
  wire  alu_io_redirect_valid; // @[EXU.scala 48:19]
  wire [63:0] alu_io_offset; // @[EXU.scala 48:19]
  wire  alu_REG_0_valid; // @[EXU.scala 48:19]
  wire [38:0] alu_REG_0_pc; // @[EXU.scala 48:19]
  wire  alu_REG_0_isMissPredict; // @[EXU.scala 48:19]
  wire [38:0] alu_REG_0_actualTarget; // @[EXU.scala 48:19]
  wire  alu_REG_0_actualTaken; // @[EXU.scala 48:19]
  wire [6:0] alu_REG_0_fuOpType; // @[EXU.scala 48:19]
  wire [1:0] alu_REG_0_btbType; // @[EXU.scala 48:19]
  wire  alu_REG_0_isRVC; // @[EXU.scala 48:19]
  wire  cnnfu_clock; // @[EXU.scala 57:21]
  wire  cnnfu_reset; // @[EXU.scala 57:21]
  wire  cnnfu_io_in_valid; // @[EXU.scala 57:21]
  wire [63:0] cnnfu_io_in_bits_src1; // @[EXU.scala 57:21]
  wire [63:0] cnnfu_io_in_bits_src2; // @[EXU.scala 57:21]
  wire [6:0] cnnfu_io_in_bits_func; // @[EXU.scala 57:21]
  wire  cnnfu_io_out_valid; // @[EXU.scala 57:21]
  wire [63:0] cnnfu_io_out_bits; // @[EXU.scala 57:21]
  wire [63:0] cnnfu_io_imm; // @[EXU.scala 57:21]
  wire [2:0] cnnfu_io_vtag; // @[EXU.scala 57:21]
  wire [3:0] cnnfu_io_length_k; // @[EXU.scala 57:21]
  wire [4:0] cnnfu_io_vec_addr; // @[EXU.scala 57:21]
  wire [1:0] cnnfu_io_algorithm; // @[EXU.scala 57:21]
  wire  cnnfu_io_loadv_valid; // @[EXU.scala 57:21]
  wire [63:0] cnnfu_io_loadv_src1; // @[EXU.scala 57:21]
  wire [63:0] cnnfu_io_loadv_src2; // @[EXU.scala 57:21]
  wire [6:0] cnnfu_io_loadv_func; // @[EXU.scala 57:21]
  wire  cnnfu_io_loadv_load_valid; // @[EXU.scala 57:21]
  wire [63:0] cnnfu_io_loadv_load_data; // @[EXU.scala 57:21]
  wire  cnnfu_io_loadv_load_exception; // @[EXU.scala 57:21]
  wire  lsu_clock; // @[EXU.scala 71:19]
  wire  lsu_reset; // @[EXU.scala 71:19]
  wire  lsu_io__in_valid; // @[EXU.scala 71:19]
  wire [63:0] lsu_io__in_bits_src1; // @[EXU.scala 71:19]
  wire [63:0] lsu_io__in_bits_src2; // @[EXU.scala 71:19]
  wire [6:0] lsu_io__in_bits_func; // @[EXU.scala 71:19]
  wire  lsu_io__out_ready; // @[EXU.scala 71:19]
  wire  lsu_io__out_valid; // @[EXU.scala 71:19]
  wire [63:0] lsu_io__out_bits; // @[EXU.scala 71:19]
  wire [63:0] lsu_io__wdata; // @[EXU.scala 71:19]
  wire [31:0] lsu_io__instr; // @[EXU.scala 71:19]
  wire  lsu_io__dmem_req_ready; // @[EXU.scala 71:19]
  wire  lsu_io__dmem_req_valid; // @[EXU.scala 71:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[EXU.scala 71:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[EXU.scala 71:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[EXU.scala 71:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[EXU.scala 71:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[EXU.scala 71:19]
  wire  lsu_io__dmem_resp_valid; // @[EXU.scala 71:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[EXU.scala 71:19]
  wire  lsu_io__dtlbPF; // @[EXU.scala 71:19]
  wire  lsu_io__loadAddrMisaligned; // @[EXU.scala 71:19]
  wire  lsu_io__storeAddrMisaligned; // @[EXU.scala 71:19]
  wire  lsu_setLr_0; // @[EXU.scala 71:19]
  wire  lsu_DTLBPF; // @[EXU.scala 71:19]
  wire  lsu_amoReq_0; // @[EXU.scala 71:19]
  wire  lsu_DTLBENABLE; // @[EXU.scala 71:19]
  wire [63:0] lsu_io_in_bits_src1; // @[EXU.scala 71:19]
  wire  lsu_DTLBFINISH; // @[EXU.scala 71:19]
  wire [63:0] lsu_setLrAddr_0; // @[EXU.scala 71:19]
  wire  lsu_setLrVal_0; // @[EXU.scala 71:19]
  wire [63:0] lsu_lr_addr; // @[EXU.scala 71:19]
  wire  mdu_clock; // @[EXU.scala 87:19]
  wire  mdu_reset; // @[EXU.scala 87:19]
  wire  mdu_io_in_ready; // @[EXU.scala 87:19]
  wire  mdu_io_in_valid; // @[EXU.scala 87:19]
  wire [63:0] mdu_io_in_bits_src1; // @[EXU.scala 87:19]
  wire [63:0] mdu_io_in_bits_src2; // @[EXU.scala 87:19]
  wire [6:0] mdu_io_in_bits_func; // @[EXU.scala 87:19]
  wire  mdu_io_out_ready; // @[EXU.scala 87:19]
  wire  mdu_io_out_valid; // @[EXU.scala 87:19]
  wire [63:0] mdu_io_out_bits; // @[EXU.scala 87:19]
  wire  csr_clock; // @[EXU.scala 92:19]
  wire  csr_reset; // @[EXU.scala 92:19]
  wire  csr_io_in_valid; // @[EXU.scala 92:19]
  wire [63:0] csr_io_in_bits_src1; // @[EXU.scala 92:19]
  wire [63:0] csr_io_in_bits_src2; // @[EXU.scala 92:19]
  wire [6:0] csr_io_in_bits_func; // @[EXU.scala 92:19]
  wire  csr_io_out_ready; // @[EXU.scala 92:19]
  wire  csr_io_out_valid; // @[EXU.scala 92:19]
  wire [63:0] csr_io_out_bits; // @[EXU.scala 92:19]
  wire [63:0] csr_io_cfIn_instr; // @[EXU.scala 92:19]
  wire [38:0] csr_io_cfIn_pc; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_0; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_1; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_2; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_3; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_4; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_5; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_6; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_7; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_8; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_9; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_10; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_intrVec_11; // @[EXU.scala 92:19]
  wire  csr_io_cfIn_crossPageIPFFix; // @[EXU.scala 92:19]
  wire [38:0] csr_io_redirect_target; // @[EXU.scala 92:19]
  wire  csr_io_redirect_valid; // @[EXU.scala 92:19]
  wire  csr_io_instrValid; // @[EXU.scala 92:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[EXU.scala 92:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 92:19]
  wire  csr_io_dmemMMU_status_sum; // @[EXU.scala 92:19]
  wire  csr_io_dmemMMU_status_mxr; // @[EXU.scala 92:19]
  wire  csr_io_dmemMMU_loadPF; // @[EXU.scala 92:19]
  wire  csr_io_dmemMMU_storePF; // @[EXU.scala 92:19]
  wire [38:0] csr_io_dmemMMU_addr; // @[EXU.scala 92:19]
  wire  csr_io_wenFix; // @[EXU.scala 92:19]
  wire  csr_set_lr; // @[EXU.scala 92:19]
  wire [63:0] csr_perfCnts_2_0; // @[EXU.scala 92:19]
  wire [63:0] csr_satp_0; // @[EXU.scala 92:19]
  wire  csr_perfCntCondMinstret; // @[EXU.scala 92:19]
  wire  csr_mtip_0; // @[EXU.scala 92:19]
  wire  csr_meip_0; // @[EXU.scala 92:19]
  wire [63:0] csr_LSUADDR; // @[EXU.scala 92:19]
  wire [11:0] csr_intrVec_0; // @[EXU.scala 92:19]
  wire  csr_msip_0; // @[EXU.scala 92:19]
  wire [63:0] csr_set_lr_addr; // @[EXU.scala 92:19]
  wire  csr_perfCntCondMultiCommit; // @[EXU.scala 92:19]
  wire  csr_set_lr_val; // @[EXU.scala 92:19]
  wire [63:0] csr_lrAddr_0; // @[EXU.scala 92:19]
  wire  mou_io_in_valid; // @[EXU.scala 106:19]
  wire [6:0] mou_io_in_bits_func; // @[EXU.scala 106:19]
  wire [38:0] mou_io_cfIn_pc; // @[EXU.scala 106:19]
  wire [38:0] mou_io_redirect_target; // @[EXU.scala 106:19]
  wire  mou_io_redirect_valid; // @[EXU.scala 106:19]
  wire  mou_flushICache_0; // @[EXU.scala 106:19]
  wire  mou_flushTLB_0; // @[EXU.scala 106:19]
  wire  _T_2 = ~io__flush; // @[EXU.scala 44:84]
  wire  fuValids_1 = io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  wire  fuValids_3 = io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  wire  fuValids_5 = io__in_bits_ctrl_fuType == 3'h5 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  wire  lsuTlbPF = lsu_io__dtlbPF;
  wire [38:0] _T_48_target = csr_io_redirect_valid ? csr_io_redirect_target : alu_io_redirect_target; // @[EXU.scala 124:10]
  wire  _T_48_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[EXU.scala 124:10]
  wire  _T_51 = 3'h1 == io__in_bits_ctrl_fuType ? lsu_io__out_valid : 1'h1; // @[Mux.scala 80:57]
  wire  _T_53 = 3'h2 == io__in_bits_ctrl_fuType ? mdu_io_out_valid : _T_51; // @[Mux.scala 80:57]
  wire  _T_55 = 3'h5 == io__in_bits_ctrl_fuType ? cnnfu_io_out_valid : _T_53; // @[Mux.scala 80:57]
  wire  _T_60 = alu_io_out_ready & alu_io_out_valid; // @[Decoupled.scala 40:37]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[ALU.scala 62:31]
  wire  _T_64 = _T_60 & ~isBru; // @[EXU.scala 152:43]
  wire  _T_66 = _T_60 & isBru; // @[EXU.scala 153:43]
  wire  _T_67 = lsu_io__out_ready & lsu_io__out_valid; // @[Decoupled.scala 40:37]
  wire  _T_68 = mdu_io_out_ready & mdu_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_69 = csr_io_out_ready & csr_io_out_valid; // @[Decoupled.scala 40:37]
  ALU alu ( // @[EXU.scala 48:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    .REG_0_valid(alu_REG_0_valid),
    .REG_0_pc(alu_REG_0_pc),
    .REG_0_isMissPredict(alu_REG_0_isMissPredict),
    .REG_0_actualTarget(alu_REG_0_actualTarget),
    .REG_0_actualTaken(alu_REG_0_actualTaken),
    .REG_0_fuOpType(alu_REG_0_fuOpType),
    .REG_0_btbType(alu_REG_0_btbType),
    .REG_0_isRVC(alu_REG_0_isRVC)
  );
  CNNFU cnnfu ( // @[EXU.scala 57:21]
    .clock(cnnfu_clock),
    .reset(cnnfu_reset),
    .io_in_valid(cnnfu_io_in_valid),
    .io_in_bits_src1(cnnfu_io_in_bits_src1),
    .io_in_bits_src2(cnnfu_io_in_bits_src2),
    .io_in_bits_func(cnnfu_io_in_bits_func),
    .io_out_valid(cnnfu_io_out_valid),
    .io_out_bits(cnnfu_io_out_bits),
    .io_imm(cnnfu_io_imm),
    .io_vtag(cnnfu_io_vtag),
    .io_length_k(cnnfu_io_length_k),
    .io_vec_addr(cnnfu_io_vec_addr),
    .io_algorithm(cnnfu_io_algorithm),
    .io_loadv_valid(cnnfu_io_loadv_valid),
    .io_loadv_src1(cnnfu_io_loadv_src1),
    .io_loadv_src2(cnnfu_io_loadv_src2),
    .io_loadv_func(cnnfu_io_loadv_func),
    .io_loadv_load_valid(cnnfu_io_loadv_load_valid),
    .io_loadv_load_data(cnnfu_io_loadv_load_data),
    .io_loadv_load_exception(cnnfu_io_loadv_load_exception)
  );
  UnpipelinedLSU lsu ( // @[EXU.scala 71:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .setLr_0(lsu_setLr_0),
    .DTLBPF(lsu_DTLBPF),
    .amoReq_0(lsu_amoReq_0),
    .DTLBENABLE(lsu_DTLBENABLE),
    .io_in_bits_src1(lsu_io_in_bits_src1),
    .DTLBFINISH(lsu_DTLBFINISH),
    .setLrAddr_0(lsu_setLrAddr_0),
    .setLrVal_0(lsu_setLrVal_0),
    .lr_addr(lsu_lr_addr)
  );
  MDU mdu ( // @[EXU.scala 87:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  CSR csr ( // @[EXU.scala 92:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_intrVec_0(csr_io_cfIn_intrVec_0),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_2(csr_io_cfIn_intrVec_2),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_4(csr_io_cfIn_intrVec_4),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_6(csr_io_cfIn_intrVec_6),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_8(csr_io_cfIn_intrVec_8),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_10(csr_io_cfIn_intrVec_10),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossPageIPFFix(csr_io_cfIn_crossPageIPFFix),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_addr(csr_io_dmemMMU_addr),
    .io_wenFix(csr_io_wenFix),
    .set_lr(csr_set_lr),
    .perfCnts_2_0(csr_perfCnts_2_0),
    .satp_0(csr_satp_0),
    .perfCntCondMinstret(csr_perfCntCondMinstret),
    .mtip_0(csr_mtip_0),
    .meip_0(csr_meip_0),
    .LSUADDR(csr_LSUADDR),
    .intrVec_0(csr_intrVec_0),
    .msip_0(csr_msip_0),
    .set_lr_addr(csr_set_lr_addr),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .set_lr_val(csr_set_lr_val),
    .lrAddr_0(csr_lrAddr_0)
  );
  MOU mou ( // @[EXU.scala 106:19]
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .flushTLB_0(mou_flushTLB_0)
  );
  assign io__in_ready = ~io__in_valid | io__out_valid; // @[EXU.scala 143:31]
  assign io__out_valid = io__in_valid & _T_55; // @[EXU.scala 130:31]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[EXU.scala 118:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target : _T_48_target; // @[EXU.scala 123:8]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid : _T_48_valid; // @[EXU.scala 123:8]
  assign io__out_bits_decode_cf_runahead_checkpoint_id = io__in_bits_cf_runahead_checkpoint_id; // @[EXU.scala 120:48]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 116:14]
  assign io__out_bits_decode_ctrl_rfWen = io__in_bits_ctrl_rfWen & (~lsuTlbPF & ~lsu_io__loadAddrMisaligned & ~
    lsu_io__storeAddrMisaligned | ~fuValids_1) & ~(csr_io_wenFix & fuValids_3); // @[EXU.scala 114:125]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 115:14]
  assign io__out_bits_commits_0 = alu_io_out_bits; // @[EXU.scala 136:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[EXU.scala 137:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[EXU.scala 139:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[EXU.scala 138:35]
  assign io__out_bits_commits_5 = cnnfu_io_out_bits; // @[EXU.scala 141:35]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[EXU.scala 78:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[EXU.scala 78:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[EXU.scala 78:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[EXU.scala 78:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[EXU.scala 78:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[EXU.scala 78:11]
  assign io__forward_valid = io__in_valid; // @[EXU.scala 145:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[EXU.scala 146:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 147:24]
  assign io__forward_wb_rfData = _T_60 ? alu_io_out_bits : lsu_io__out_bits; // @[EXU.scala 148:30]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 149:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[EXU.scala 103:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 104:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[EXU.scala 104:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[EXU.scala 104:18]
  assign flushICache = mou_flushICache_0;
  assign perfCnts_2 = csr_perfCnts_2_0;
  assign satp = csr_satp_0;
  assign REG_0_valid = alu_REG_0_valid;
  assign REG_0_pc = alu_REG_0_pc;
  assign REG_0_isMissPredict = alu_REG_0_isMissPredict;
  assign REG_0_actualTarget = alu_REG_0_actualTarget;
  assign REG_0_actualTaken = alu_REG_0_actualTaken;
  assign REG_0_fuOpType = alu_REG_0_fuOpType;
  assign REG_0_btbType = alu_REG_0_btbType;
  assign REG_0_isRVC = alu_REG_0_isRVC;
  assign amoReq = lsu_amoReq_0;
  assign intrVec = csr_intrVec_0;
  assign flushTLB = mou_flushTLB_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = io__in_bits_ctrl_fuType == 3'h0 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  assign alu_io_in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 38:34]
  assign alu_io_in_bits_src2 = io__in_bits_data_src2; // @[EXU.scala 39:34]
  assign alu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[ALU.scala 83:15]
  assign alu_io_out_ready = 1'h1; // @[EXU.scala 52:20]
  assign alu_io_cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 50:15]
  assign alu_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 50:15]
  assign alu_io_cfIn_pnpc = io__in_bits_cf_pnpc; // @[EXU.scala 50:15]
  assign alu_io_cfIn_brIdx = io__in_bits_cf_brIdx; // @[EXU.scala 50:15]
  assign alu_io_offset = io__in_bits_data_imm; // @[EXU.scala 51:17]
  assign cnnfu_clock = clock;
  assign cnnfu_reset = reset;
  assign cnnfu_io_in_valid = io__in_bits_ctrl_fuType == 3'h5 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  assign cnnfu_io_in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 38:34]
  assign cnnfu_io_in_bits_src2 = io__in_bits_data_src2; // @[EXU.scala 39:34]
  assign cnnfu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[CNN_FU.scala 70:15]
  assign cnnfu_io_imm = io__in_bits_data_imm; // @[EXU.scala 59:16]
  assign cnnfu_io_vtag = io__in_bits_ctrl_vtag; // @[EXU.scala 60:17]
  assign cnnfu_io_length_k = io__in_bits_ctrl_length_k; // @[EXU.scala 62:21]
  assign cnnfu_io_vec_addr = io__in_bits_ctrl_vec_addr; // @[EXU.scala 61:21]
  assign cnnfu_io_algorithm = io__in_bits_ctrl_algorithm; // @[EXU.scala 63:22]
  assign cnnfu_io_loadv_load_valid = lsu_io__out_valid; // @[EXU.scala 82:29]
  assign cnnfu_io_loadv_load_data = lsu_io__out_bits; // @[EXU.scala 83:28]
  assign cnnfu_io_loadv_load_exception = lsuTlbPF | lsu_io__loadAddrMisaligned | lsu_io__storeAddrMisaligned; // @[EXU.scala 84:74]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = fuValids_5 ? cnnfu_io_loadv_valid : fuValids_1; // @[EXU.scala 66:22]
  assign lsu_io__in_bits_src1 = fuValids_5 ? cnnfu_io_loadv_src1 : io__in_bits_data_src1; // @[EXU.scala 67:21]
  assign lsu_io__in_bits_src2 = fuValids_5 ? cnnfu_io_loadv_src2 : io__in_bits_data_imm; // @[EXU.scala 68:21]
  assign lsu_io__in_bits_func = fuValids_5 ? cnnfu_io_loadv_func : io__in_bits_ctrl_fuOpType; // @[EXU.scala 69:21]
  assign lsu_io__out_ready = 1'h1; // @[EXU.scala 79:20]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[EXU.scala 39:34]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[EXU.scala 76:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[EXU.scala 78:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[EXU.scala 78:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[EXU.scala 78:11]
  assign lsu_DTLBPF = _T_28_0;
  assign lsu_DTLBENABLE = vmEnable;
  assign lsu_DTLBFINISH = _T_27_0;
  assign lsu_lr_addr = csr_lrAddr_0;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = io__in_bits_ctrl_fuType == 3'h2 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 38:34]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[EXU.scala 39:34]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[EXU.scala 89:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 38:34]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[EXU.scala 39:34]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[CSR.scala 200:15]
  assign csr_io_out_ready = 1'h1; // @[EXU.scala 101:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 94:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 94:15]
  assign csr_io_cfIn_exceptionVec_1 = io__in_bits_cf_exceptionVec_1; // @[EXU.scala 94:15]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[EXU.scala 94:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[EXU.scala 95:48]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[EXU.scala 96:49]
  assign csr_io_cfIn_exceptionVec_12 = io__in_bits_cf_exceptionVec_12; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_0 = io__in_bits_cf_intrVec_0; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_2 = io__in_bits_cf_intrVec_2; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_4 = io__in_bits_cf_intrVec_4; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_6 = io__in_bits_cf_intrVec_6; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_8 = io__in_bits_cf_intrVec_8; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_10 = io__in_bits_cf_intrVec_10; // @[EXU.scala 94:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[EXU.scala 94:15]
  assign csr_io_cfIn_crossPageIPFFix = io__in_bits_cf_crossPageIPFFix; // @[EXU.scala 94:15]
  assign csr_io_instrValid = io__in_valid & _T_2; // @[EXU.scala 97:36]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[EXU.scala 104:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[EXU.scala 104:18]
  assign csr_io_dmemMMU_addr = io__memMMU_dmem_addr; // @[EXU.scala 104:18]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_LSUADDR = lsu_io_in_bits_src1;
  assign csr_msip_0 = io_extra_msip;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign mou_io_in_valid = io__in_bits_ctrl_fuType == 3'h4 & io__in_valid & ~io__flush; // @[EXU.scala 44:81]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 109:15]
endmodule
module WBU(
  input         clock,
  input         io__in_valid,
  input  [38:0] io__in_bits_decode_cf_pc,
  input  [38:0] io__in_bits_decode_cf_redirect_target,
  input         io__in_bits_decode_cf_redirect_valid,
  input  [63:0] io__in_bits_decode_cf_runahead_checkpoint_id,
  input  [2:0]  io__in_bits_decode_ctrl_fuType,
  input         io__in_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_bits_decode_ctrl_rfDest,
  input  [63:0] io__in_bits_commits_0,
  input  [63:0] io__in_bits_commits_1,
  input  [63:0] io__in_bits_commits_2,
  input  [63:0] io__in_bits_commits_3,
  input  [63:0] io__in_bits_commits_5,
  output        io__wb_rfWen,
  output [4:0]  io__wb_rfDest,
  output [63:0] io__wb_rfData,
  output [38:0] io__redirect_target,
  output        io__redirect_valid,
  output [38:0] io_in_bits_decode_cf_pc,
  output [4:0]  io_wb_rfDest,
  output        io_in_valid,
  output        io_wb_rfWen,
  output [63:0] io_wb_rfData,
  output        io_in_valid_0,
  output        falseWire_0
);
  wire  runahead_redirect_io_clock; // @[WBU.scala 41:33]
  wire [7:0] runahead_redirect_io_coreid; // @[WBU.scala 41:33]
  wire  runahead_redirect_io_valid; // @[WBU.scala 41:33]
  wire [63:0] runahead_redirect_io_pc; // @[WBU.scala 41:33]
  wire [63:0] runahead_redirect_io_target_pc; // @[WBU.scala 41:33]
  wire [63:0] runahead_redirect_io_checkpoint_id; // @[WBU.scala 41:33]
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[WBU.scala 34:{16,16}]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[WBU.scala 34:{16,16}]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[WBU.scala 34:{16,16}]
  wire [63:0] _GEN_4 = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[WBU.scala 34:{16,16}]
  wire  falseWire = 1'h0;
  DifftestRunaheadRedirectEvent runahead_redirect ( // @[WBU.scala 41:33]
    .io_clock(runahead_redirect_io_clock),
    .io_coreid(runahead_redirect_io_coreid),
    .io_valid(runahead_redirect_io_valid),
    .io_pc(runahead_redirect_io_pc),
    .io_target_pc(runahead_redirect_io_target_pc),
    .io_checkpoint_id(runahead_redirect_io_checkpoint_id)
  );
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[WBU.scala 32:47]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[WBU.scala 33:16]
  assign io__wb_rfData = 3'h5 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_5 : _GEN_4; // @[WBU.scala 34:{16,16}]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[WBU.scala 38:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[WBU.scala 39:60]
  assign io_in_bits_decode_cf_pc = io__in_bits_decode_cf_pc;
  assign io_wb_rfDest = io__wb_rfDest;
  assign io_in_valid = io__in_valid;
  assign io_wb_rfWen = io__wb_rfWen;
  assign io_wb_rfData = io__wb_rfData;
  assign io_in_valid_0 = io__in_valid;
  assign falseWire_0 = falseWire;
  assign runahead_redirect_io_clock = clock; // @[WBU.scala 42:30]
  assign runahead_redirect_io_coreid = 8'h0; // @[WBU.scala 43:31]
  assign runahead_redirect_io_valid = io__redirect_valid; // @[WBU.scala 44:30]
  assign runahead_redirect_io_pc = {{25'd0}, io__in_bits_decode_cf_pc}; // @[WBU.scala 45:27]
  assign runahead_redirect_io_target_pc = {{25'd0}, io__in_bits_decode_cf_redirect_target}; // @[WBU.scala 46:34]
  assign runahead_redirect_io_checkpoint_id = io__in_bits_decode_cf_runahead_checkpoint_id; // @[WBU.scala 47:38]
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input  [63:0] io_in_0_bits_cf_runahead_checkpoint_id,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input  [2:0]  io_in_0_bits_ctrl_vtag,
  input  [4:0]  io_in_0_bits_ctrl_vec_addr,
  input  [3:0]  io_in_0_bits_ctrl_length_k,
  input  [1:0]  io_in_0_bits_ctrl_algorithm,
  input  [63:0] io_in_0_bits_data_imm,
  input  [1:0]  io_flush,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  output [1:0]  io_memMMU_imem_priviledgeMode,
  output [1:0]  io_memMMU_dmem_priviledgeMode,
  output        io_memMMU_dmem_status_sum,
  output        io_memMMU_dmem_status_mxr,
  input         io_memMMU_dmem_loadPF,
  input         io_memMMU_dmem_storePF,
  input  [38:0] io_memMMU_dmem_addr,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         _T_28,
  output        flushICache,
  output [63:0] perfCnts_2,
  output [38:0] io_in_bits_decode_cf_pc,
  output [63:0] satp,
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output        REG_0_actualTaken,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC,
  output [4:0]  io_wb_rfDest,
  input         io_extra_mtip,
  output        amoReq,
  input         io_extra_meip_0,
  input         vmEnable,
  output        io_wb_rfWen,
  output [63:0] io_wb_rfData,
  output [11:0] intrVec,
  input         _T_27,
  input         io_extra_msip,
  output        flushTLB,
  output        io_in_valid_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[Backend.scala 680:20]
  wire  isu_reset; // @[Backend.scala 680:20]
  wire  isu_io_in_0_ready; // @[Backend.scala 680:20]
  wire  isu_io_in_0_valid; // @[Backend.scala 680:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[Backend.scala 680:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[Backend.scala 680:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_0; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_2; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_4; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_6; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_8; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_10; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[Backend.scala 680:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 680:20]
  wire [63:0] isu_io_in_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[Backend.scala 680:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[Backend.scala 680:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 680:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 680:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 680:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[Backend.scala 680:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[Backend.scala 680:20]
  wire [2:0] isu_io_in_0_bits_ctrl_vtag; // @[Backend.scala 680:20]
  wire [4:0] isu_io_in_0_bits_ctrl_vec_addr; // @[Backend.scala 680:20]
  wire [3:0] isu_io_in_0_bits_ctrl_length_k; // @[Backend.scala 680:20]
  wire [1:0] isu_io_in_0_bits_ctrl_algorithm; // @[Backend.scala 680:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[Backend.scala 680:20]
  wire  isu_io_out_ready; // @[Backend.scala 680:20]
  wire  isu_io_out_valid; // @[Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[Backend.scala 680:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[Backend.scala 680:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_0; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_2; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_4; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_6; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_8; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_10; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[Backend.scala 680:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_cf_crossPageIPFFix; // @[Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_cf_runahead_checkpoint_id; // @[Backend.scala 680:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[Backend.scala 680:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[Backend.scala 680:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[Backend.scala 680:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[Backend.scala 680:20]
  wire [2:0] isu_io_out_bits_ctrl_vtag; // @[Backend.scala 680:20]
  wire [4:0] isu_io_out_bits_ctrl_vec_addr; // @[Backend.scala 680:20]
  wire [3:0] isu_io_out_bits_ctrl_length_k; // @[Backend.scala 680:20]
  wire [1:0] isu_io_out_bits_ctrl_algorithm; // @[Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[Backend.scala 680:20]
  wire  isu_io_wb_rfWen; // @[Backend.scala 680:20]
  wire [4:0] isu_io_wb_rfDest; // @[Backend.scala 680:20]
  wire [63:0] isu_io_wb_rfData; // @[Backend.scala 680:20]
  wire  isu_io_forward_valid; // @[Backend.scala 680:20]
  wire  isu_io_forward_wb_rfWen; // @[Backend.scala 680:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[Backend.scala 680:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[Backend.scala 680:20]
  wire [2:0] isu_io_forward_fuType; // @[Backend.scala 680:20]
  wire  isu_io_flush; // @[Backend.scala 680:20]
  wire  exu_clock; // @[Backend.scala 681:20]
  wire  exu_reset; // @[Backend.scala 681:20]
  wire  exu_io__in_ready; // @[Backend.scala 681:20]
  wire  exu_io__in_valid; // @[Backend.scala 681:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[Backend.scala 681:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[Backend.scala 681:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_0; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_2; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_4; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_6; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_8; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_10; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[Backend.scala 681:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_cf_crossPageIPFFix; // @[Backend.scala 681:20]
  wire [63:0] exu_io__in_bits_cf_runahead_checkpoint_id; // @[Backend.scala 681:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[Backend.scala 681:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[Backend.scala 681:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[Backend.scala 681:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[Backend.scala 681:20]
  wire [2:0] exu_io__in_bits_ctrl_vtag; // @[Backend.scala 681:20]
  wire [4:0] exu_io__in_bits_ctrl_vec_addr; // @[Backend.scala 681:20]
  wire [3:0] exu_io__in_bits_ctrl_length_k; // @[Backend.scala 681:20]
  wire [1:0] exu_io__in_bits_ctrl_algorithm; // @[Backend.scala 681:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[Backend.scala 681:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[Backend.scala 681:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[Backend.scala 681:20]
  wire  exu_io__out_ready; // @[Backend.scala 681:20]
  wire  exu_io__out_valid; // @[Backend.scala 681:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[Backend.scala 681:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[Backend.scala 681:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[Backend.scala 681:20]
  wire [63:0] exu_io__out_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 681:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[Backend.scala 681:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[Backend.scala 681:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[Backend.scala 681:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[Backend.scala 681:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[Backend.scala 681:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[Backend.scala 681:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[Backend.scala 681:20]
  wire [63:0] exu_io__out_bits_commits_5; // @[Backend.scala 681:20]
  wire  exu_io__flush; // @[Backend.scala 681:20]
  wire  exu_io__dmem_req_ready; // @[Backend.scala 681:20]
  wire  exu_io__dmem_req_valid; // @[Backend.scala 681:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[Backend.scala 681:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[Backend.scala 681:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[Backend.scala 681:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[Backend.scala 681:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[Backend.scala 681:20]
  wire  exu_io__dmem_resp_valid; // @[Backend.scala 681:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[Backend.scala 681:20]
  wire  exu_io__forward_valid; // @[Backend.scala 681:20]
  wire  exu_io__forward_wb_rfWen; // @[Backend.scala 681:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[Backend.scala 681:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[Backend.scala 681:20]
  wire [2:0] exu_io__forward_fuType; // @[Backend.scala 681:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 681:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 681:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[Backend.scala 681:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 681:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[Backend.scala 681:20]
  wire  exu_io__memMMU_dmem_storePF; // @[Backend.scala 681:20]
  wire [38:0] exu_io__memMMU_dmem_addr; // @[Backend.scala 681:20]
  wire  exu__T_28_0; // @[Backend.scala 681:20]
  wire  exu_flushICache; // @[Backend.scala 681:20]
  wire [63:0] exu_perfCnts_2; // @[Backend.scala 681:20]
  wire [63:0] exu_satp; // @[Backend.scala 681:20]
  wire  exu_REG_0_valid; // @[Backend.scala 681:20]
  wire [38:0] exu_REG_0_pc; // @[Backend.scala 681:20]
  wire  exu_REG_0_isMissPredict; // @[Backend.scala 681:20]
  wire [38:0] exu_REG_0_actualTarget; // @[Backend.scala 681:20]
  wire  exu_REG_0_actualTaken; // @[Backend.scala 681:20]
  wire [6:0] exu_REG_0_fuOpType; // @[Backend.scala 681:20]
  wire [1:0] exu_REG_0_btbType; // @[Backend.scala 681:20]
  wire  exu_REG_0_isRVC; // @[Backend.scala 681:20]
  wire  exu_io_in_valid; // @[Backend.scala 681:20]
  wire  exu_io_extra_mtip; // @[Backend.scala 681:20]
  wire  exu_amoReq; // @[Backend.scala 681:20]
  wire  exu_io_extra_meip_0; // @[Backend.scala 681:20]
  wire  exu_vmEnable; // @[Backend.scala 681:20]
  wire [11:0] exu_intrVec; // @[Backend.scala 681:20]
  wire  exu__T_27_0; // @[Backend.scala 681:20]
  wire  exu_io_extra_msip; // @[Backend.scala 681:20]
  wire  exu_flushTLB; // @[Backend.scala 681:20]
  wire  exu_falseWire; // @[Backend.scala 681:20]
  wire  wbu_clock; // @[Backend.scala 682:20]
  wire  wbu_io__in_valid; // @[Backend.scala 682:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[Backend.scala 682:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[Backend.scala 682:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_decode_cf_runahead_checkpoint_id; // @[Backend.scala 682:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[Backend.scala 682:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[Backend.scala 682:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_5; // @[Backend.scala 682:20]
  wire  wbu_io__wb_rfWen; // @[Backend.scala 682:20]
  wire [4:0] wbu_io__wb_rfDest; // @[Backend.scala 682:20]
  wire [63:0] wbu_io__wb_rfData; // @[Backend.scala 682:20]
  wire [38:0] wbu_io__redirect_target; // @[Backend.scala 682:20]
  wire  wbu_io__redirect_valid; // @[Backend.scala 682:20]
  wire [38:0] wbu_io_in_bits_decode_cf_pc; // @[Backend.scala 682:20]
  wire [4:0] wbu_io_wb_rfDest; // @[Backend.scala 682:20]
  wire  wbu_io_in_valid; // @[Backend.scala 682:20]
  wire  wbu_io_wb_rfWen; // @[Backend.scala 682:20]
  wire [63:0] wbu_io_wb_rfData; // @[Backend.scala 682:20]
  wire  wbu_io_in_valid_0; // @[Backend.scala 682:20]
  wire  wbu_falseWire_0; // @[Backend.scala 682:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = isu_io_out_valid & exu_io__in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = isu_io_out_valid & exu_io__in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [63:0] r_cf_instr; // @[Reg.scala 15:16]
  reg [38:0] r_cf_pc; // @[Reg.scala 15:16]
  reg [38:0] r_cf_pnpc; // @[Reg.scala 15:16]
  reg  r_cf_exceptionVec_1; // @[Reg.scala 15:16]
  reg  r_cf_exceptionVec_2; // @[Reg.scala 15:16]
  reg  r_cf_exceptionVec_12; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_0; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_1; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_2; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_3; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_4; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_5; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_6; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_7; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_8; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_9; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_10; // @[Reg.scala 15:16]
  reg  r_cf_intrVec_11; // @[Reg.scala 15:16]
  reg [3:0] r_cf_brIdx; // @[Reg.scala 15:16]
  reg  r_cf_crossPageIPFFix; // @[Reg.scala 15:16]
  reg [63:0] r_cf_runahead_checkpoint_id; // @[Reg.scala 15:16]
  reg [2:0] r_ctrl_fuType; // @[Reg.scala 15:16]
  reg [6:0] r_ctrl_fuOpType; // @[Reg.scala 15:16]
  reg  r_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] r_ctrl_rfDest; // @[Reg.scala 15:16]
  reg [2:0] r_ctrl_vtag; // @[Reg.scala 15:16]
  reg [4:0] r_ctrl_vec_addr; // @[Reg.scala 15:16]
  reg [3:0] r_ctrl_length_k; // @[Reg.scala 15:16]
  reg [1:0] r_ctrl_algorithm; // @[Reg.scala 15:16]
  reg [63:0] r_data_src1; // @[Reg.scala 15:16]
  reg [63:0] r_data_src2; // @[Reg.scala 15:16]
  reg [63:0] r_data_imm; // @[Reg.scala 15:16]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _T_5 = exu_io__out_valid; // @[Pipeline.scala 26:22]
  reg [38:0] r_1_decode_cf_pc; // @[Reg.scala 15:16]
  reg [38:0] r_1_decode_cf_redirect_target; // @[Reg.scala 15:16]
  reg  r_1_decode_cf_redirect_valid; // @[Reg.scala 15:16]
  reg [63:0] r_1_decode_cf_runahead_checkpoint_id; // @[Reg.scala 15:16]
  reg [2:0] r_1_decode_ctrl_fuType; // @[Reg.scala 15:16]
  reg  r_1_decode_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] r_1_decode_ctrl_rfDest; // @[Reg.scala 15:16]
  reg [63:0] r_1_commits_0; // @[Reg.scala 15:16]
  reg [63:0] r_1_commits_1; // @[Reg.scala 15:16]
  reg [63:0] r_1_commits_2; // @[Reg.scala 15:16]
  reg [63:0] r_1_commits_3; // @[Reg.scala 15:16]
  reg [63:0] r_1_commits_5; // @[Reg.scala 15:16]
  ISU isu ( // @[Backend.scala 680:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(isu_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(isu_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(isu_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(isu_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(isu_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(isu_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(isu_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_cf_runahead_checkpoint_id(isu_io_in_0_bits_cf_runahead_checkpoint_id),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_vtag(isu_io_in_0_bits_ctrl_vtag),
    .io_in_0_bits_ctrl_vec_addr(isu_io_in_0_bits_ctrl_vec_addr),
    .io_in_0_bits_ctrl_length_k(isu_io_in_0_bits_ctrl_length_k),
    .io_in_0_bits_ctrl_algorithm(isu_io_in_0_bits_ctrl_algorithm),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(isu_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(isu_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(isu_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(isu_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(isu_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(isu_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(isu_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_cf_runahead_checkpoint_id(isu_io_out_bits_cf_runahead_checkpoint_id),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_vtag(isu_io_out_bits_ctrl_vtag),
    .io_out_bits_ctrl_vec_addr(isu_io_out_bits_ctrl_vec_addr),
    .io_out_bits_ctrl_length_k(isu_io_out_bits_ctrl_length_k),
    .io_out_bits_ctrl_algorithm(isu_io_out_bits_ctrl_algorithm),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush)
  );
  EXU exu ( // @[Backend.scala 681:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_0(exu_io__in_bits_cf_intrVec_0),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_2(exu_io__in_bits_cf_intrVec_2),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_4(exu_io__in_bits_cf_intrVec_4),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_6(exu_io__in_bits_cf_intrVec_6),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_8(exu_io__in_bits_cf_intrVec_8),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_10(exu_io__in_bits_cf_intrVec_10),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossPageIPFFix(exu_io__in_bits_cf_crossPageIPFFix),
    .io__in_bits_cf_runahead_checkpoint_id(exu_io__in_bits_cf_runahead_checkpoint_id),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_ctrl_vtag(exu_io__in_bits_ctrl_vtag),
    .io__in_bits_ctrl_vec_addr(exu_io__in_bits_ctrl_vec_addr),
    .io__in_bits_ctrl_length_k(exu_io__in_bits_ctrl_length_k),
    .io__in_bits_ctrl_algorithm(exu_io__in_bits_ctrl_algorithm),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_cf_runahead_checkpoint_id(exu_io__out_bits_decode_cf_runahead_checkpoint_id),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__out_bits_commits_5(exu_io__out_bits_commits_5),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_addr(exu_io__memMMU_dmem_addr),
    ._T_28_0(exu__T_28_0),
    .flushICache(exu_flushICache),
    .perfCnts_2(exu_perfCnts_2),
    .satp(exu_satp),
    .REG_0_valid(exu_REG_0_valid),
    .REG_0_pc(exu_REG_0_pc),
    .REG_0_isMissPredict(exu_REG_0_isMissPredict),
    .REG_0_actualTarget(exu_REG_0_actualTarget),
    .REG_0_actualTaken(exu_REG_0_actualTaken),
    .REG_0_fuOpType(exu_REG_0_fuOpType),
    .REG_0_btbType(exu_REG_0_btbType),
    .REG_0_isRVC(exu_REG_0_isRVC),
    .io_in_valid(exu_io_in_valid),
    .io_extra_mtip(exu_io_extra_mtip),
    .amoReq(exu_amoReq),
    .io_extra_meip_0(exu_io_extra_meip_0),
    .vmEnable(exu_vmEnable),
    .intrVec(exu_intrVec),
    ._T_27_0(exu__T_27_0),
    .io_extra_msip(exu_io_extra_msip),
    .flushTLB(exu_flushTLB),
    .falseWire(exu_falseWire)
  );
  WBU wbu ( // @[Backend.scala 682:20]
    .clock(wbu_clock),
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_cf_runahead_checkpoint_id(wbu_io__in_bits_decode_cf_runahead_checkpoint_id),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__in_bits_commits_5(wbu_io__in_bits_commits_5),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .io_in_bits_decode_cf_pc(wbu_io_in_bits_decode_cf_pc),
    .io_wb_rfDest(wbu_io_wb_rfDest),
    .io_in_valid(wbu_io_in_valid),
    .io_wb_rfWen(wbu_io_wb_rfWen),
    .io_wb_rfData(wbu_io_wb_rfData),
    .io_in_valid_0(wbu_io_in_valid_0),
    .falseWire_0(wbu_falseWire_0)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[Backend.scala 687:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[Backend.scala 699:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[Backend.scala 699:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[Backend.scala 699:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[Backend.scala 699:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[Backend.scala 699:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[Backend.scala 699:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 697:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 698:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[Backend.scala 698:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 698:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[Backend.scala 693:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[Backend.scala 693:15]
  assign flushICache = exu_flushICache;
  assign perfCnts_2 = exu_perfCnts_2;
  assign io_in_bits_decode_cf_pc = wbu_io_in_bits_decode_cf_pc;
  assign satp = exu_satp;
  assign REG_0_valid = exu_REG_0_valid;
  assign REG_0_pc = exu_REG_0_pc;
  assign REG_0_isMissPredict = exu_REG_0_isMissPredict;
  assign REG_0_actualTarget = exu_REG_0_actualTarget;
  assign REG_0_actualTaken = exu_REG_0_actualTaken;
  assign REG_0_fuOpType = exu_REG_0_fuOpType;
  assign REG_0_btbType = exu_REG_0_btbType;
  assign REG_0_isRVC = exu_REG_0_isRVC;
  assign io_wb_rfDest = wbu_io_wb_rfDest;
  assign amoReq = exu_amoReq;
  assign io_wb_rfWen = wbu_io_wb_rfWen;
  assign io_wb_rfData = wbu_io_wb_rfData;
  assign intrVec = exu_intrVec;
  assign flushTLB = exu_flushTLB;
  assign io_in_valid_0 = wbu_io_in_valid_0;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_runahead_checkpoint_id = io_in_0_bits_cf_runahead_checkpoint_id; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_vtag = io_in_0_bits_ctrl_vtag; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_vec_addr = io_in_0_bits_ctrl_vec_addr; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_length_k = io_in_0_bits_ctrl_length_k; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_algorithm = io_in_0_bits_ctrl_algorithm; // @[Backend.scala 687:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[Backend.scala 687:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[Backend.scala 692:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[Backend.scala 692:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[Backend.scala 692:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[Backend.scala 695:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[Backend.scala 695:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[Backend.scala 695:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[Backend.scala 695:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[Backend.scala 695:18]
  assign isu_io_flush = io_flush[0]; // @[Backend.scala 689:27]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = REG; // @[Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = r_cf_instr; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = r_cf_pc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = r_cf_pnpc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = r_cf_exceptionVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = r_cf_exceptionVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = r_cf_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_0 = r_cf_intrVec_0; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = r_cf_intrVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_2 = r_cf_intrVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = r_cf_intrVec_3; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_4 = r_cf_intrVec_4; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = r_cf_intrVec_5; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_6 = r_cf_intrVec_6; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = r_cf_intrVec_7; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_8 = r_cf_intrVec_8; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = r_cf_intrVec_9; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_10 = r_cf_intrVec_10; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = r_cf_intrVec_11; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = r_cf_brIdx; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossPageIPFFix = r_cf_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_runahead_checkpoint_id = r_cf_runahead_checkpoint_id; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = r_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = r_ctrl_fuOpType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = r_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = r_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_vtag = r_ctrl_vtag; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_vec_addr = r_ctrl_vec_addr; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_length_k = r_ctrl_length_k; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_algorithm = r_ctrl_algorithm; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = r_data_src1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = r_data_src2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = r_data_imm; // @[Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[Backend.scala 690:27]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[Backend.scala 699:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[Backend.scala 699:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[Backend.scala 699:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[Backend.scala 698:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[Backend.scala 698:18]
  assign exu_io__memMMU_dmem_addr = io_memMMU_dmem_addr; // @[Backend.scala 698:18]
  assign exu__T_28_0 = _T_28;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu_vmEnable = vmEnable;
  assign exu__T_27_0 = _T_27;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu_falseWire = wbu_falseWire_0;
  assign wbu_clock = clock;
  assign wbu_io__in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_pc = r_1_decode_cf_pc; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = r_1_decode_cf_redirect_target; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = r_1_decode_cf_redirect_valid; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_runahead_checkpoint_id = r_1_decode_cf_runahead_checkpoint_id; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = r_1_decode_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = r_1_decode_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = r_1_decode_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = r_1_commits_0; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = r_1_commits_1; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = r_1_commits_2; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = r_1_commits_3; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_5 = r_1_commits_5; // @[Pipeline.scala 30:16]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_instr <= isu_io_out_bits_cf_instr; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_pc <= isu_io_out_bits_cf_pc; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_pnpc <= isu_io_out_bits_cf_pnpc; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_0 <= isu_io_out_bits_cf_intrVec_0; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_2 <= isu_io_out_bits_cf_intrVec_2; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_4 <= isu_io_out_bits_cf_intrVec_4; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_6 <= isu_io_out_bits_cf_intrVec_6; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_8 <= isu_io_out_bits_cf_intrVec_8; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_10 <= isu_io_out_bits_cf_intrVec_10; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_brIdx <= isu_io_out_bits_cf_brIdx; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_crossPageIPFFix <= isu_io_out_bits_cf_crossPageIPFFix; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_cf_runahead_checkpoint_id <= isu_io_out_bits_cf_runahead_checkpoint_id; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_fuType <= isu_io_out_bits_ctrl_fuType; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_vtag <= isu_io_out_bits_ctrl_vtag; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_vec_addr <= isu_io_out_bits_ctrl_vec_addr; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_length_k <= isu_io_out_bits_ctrl_length_k; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_ctrl_algorithm <= isu_io_out_bits_ctrl_algorithm; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_data_src1 <= isu_io_out_bits_data_src1; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_data_src2 <= isu_io_out_bits_data_src2; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_data_imm <= isu_io_out_bits_data_imm; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[Pipeline.scala 27:20]
      REG_1 <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG_1 <= _T_5;
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_decode_cf_pc <= exu_io__out_bits_decode_cf_pc; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_decode_cf_runahead_checkpoint_id <= exu_io__out_bits_decode_cf_runahead_checkpoint_id; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_commits_0 <= exu_io__out_bits_commits_0; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_commits_1 <= exu_io__out_bits_commits_1; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_commits_2 <= exu_io__out_bits_commits_2; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_commits_3 <= exu_io__out_bits_commits_3; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_commits_5 <= exu_io__out_bits_commits_5; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  r_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  r_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_cf_exceptionVec_12 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_cf_intrVec_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_cf_intrVec_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_cf_intrVec_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_cf_intrVec_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_cf_intrVec_4 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_cf_intrVec_5 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_cf_intrVec_6 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_cf_intrVec_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_cf_intrVec_8 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_cf_intrVec_9 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_cf_intrVec_10 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_cf_intrVec_11 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_cf_brIdx = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  r_cf_crossPageIPFFix = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  r_cf_runahead_checkpoint_id = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  r_ctrl_fuType = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  r_ctrl_fuOpType = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  r_ctrl_rfWen = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_ctrl_rfDest = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  r_ctrl_vtag = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  r_ctrl_vec_addr = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  r_ctrl_length_k = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  r_ctrl_algorithm = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  r_data_src1 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  r_data_src2 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  r_data_imm = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  REG_1 = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  r_1_decode_cf_pc = _RAND_34[38:0];
  _RAND_35 = {2{`RANDOM}};
  r_1_decode_cf_redirect_target = _RAND_35[38:0];
  _RAND_36 = {1{`RANDOM}};
  r_1_decode_cf_redirect_valid = _RAND_36[0:0];
  _RAND_37 = {2{`RANDOM}};
  r_1_decode_cf_runahead_checkpoint_id = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  r_1_decode_ctrl_fuType = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  r_1_decode_ctrl_rfWen = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_1_decode_ctrl_rfDest = _RAND_40[4:0];
  _RAND_41 = {2{`RANDOM}};
  r_1_commits_0 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  r_1_commits_1 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  r_1_commits_2 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  r_1_commits_3 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  r_1_commits_5 = _RAND_45[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] value; // @[Counter.scala 60:40]
  reg  lockIdx; // @[Arbiter.scala 46:22]
  wire  locked = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire  choice = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 88:{27,36}]
  wire  _T_2 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[Arbiter.scala 57:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : io_in_0_bits_wmask; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:{15,15}]
  assign io_chosen = locked ? lockIdx : choice; // @[Arbiter.scala 40:13 55:{19,31}]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      lockIdx <= io_chosen; // @[Arbiter.scala 51:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [3:0]  io_in_0_resp_bits_cmd,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [2:0]  io_in_1_req_bits_size,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [7:0]  io_in_1_req_bits_wmask,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [3:0]  io_in_1_resp_bits_cmd,
  output [63:0] io_in_1_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  reg  inflightSrc; // @[Crossbar.scala 105:24]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_25 | _T_26 ? 2'h2 : state; // @[Crossbar.scala 124:{80,88} 98:22]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [1:0] _GEN_9 = _T_29 ? 2'h0 : state; // @[Crossbar.scala 128:{50,58} 98:22]
  LockingArbiter inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:{13,13} 113:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:{13,13} 113:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[Crossbar.scala 109:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = 1'h1; // @[Crossbar.scala 116:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:37]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 98:22]
      state <= 2'h0; // @[Crossbar.scala 98:22]
    end else if (2'h0 == state) begin // @[Crossbar.scala 119:18]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        if (_T_4) begin // @[Crossbar.scala 123:38]
          state <= 2'h1; // @[Crossbar.scala 123:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (2'h1 == state) begin // @[Crossbar.scala 119:18]
      if (_T_29 & _T_30) begin // @[Crossbar.scala 127:82]
        state <= 2'h0; // @[Crossbar.scala 127:90]
      end
    end else if (2'h2 == state) begin // @[Crossbar.scala 119:18]
      state <= _GEN_9;
    end
    if (2'h0 == state) begin // @[Crossbar.scala 119:18]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        inflightSrc <= inputArb_io_chosen; // @[Crossbar.scala 122:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [3:0]  io_in_1_bits_cmd,
  input  [63:0] io_in_1_bits_wdata,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [3:0]  io_in_2_bits_cmd,
  input  [63:0] io_in_2_bits_wdata,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input  [2:0]  io_in_3_bits_size,
  input  [3:0]  io_in_3_bits_cmd,
  input  [7:0]  io_in_3_bits_wmask,
  input  [63:0] io_in_3_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 41:{16,16}]
  wire [63:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:{15,15}]
  wire [63:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_5; // @[Arbiter.scala 42:{15,15}]
  wire [7:0] _GEN_9 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[Arbiter.scala 42:{15,15}]
  wire [7:0] _GEN_10 = 2'h2 == io_chosen ? 8'hff : _GEN_9; // @[Arbiter.scala 42:{15,15}]
  wire [3:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:{15,15}]
  wire [3:0] _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_13; // @[Arbiter.scala 42:{15,15}]
  wire [2:0] _GEN_17 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[Arbiter.scala 42:{15,15}]
  wire [2:0] _GEN_18 = 2'h2 == io_chosen ? 3'h3 : _GEN_17; // @[Arbiter.scala 42:{15,15}]
  wire [31:0] _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:{15,15}]
  wire [31:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_21; // @[Arbiter.scala 42:{15,15}]
  reg [2:0] value; // @[Counter.scala 60:40]
  reg [1:0] lockIdx; // @[Arbiter.scala 46:22]
  wire  locked = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [1:0] _GEN_27 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 88:{27,36}]
  wire [1:0] _GEN_28 = io_in_1_valid ? 2'h1 : _GEN_27; // @[Arbiter.scala 88:{27,36}]
  wire [1:0] choice = io_in_0_valid ? 2'h0 : _GEN_28; // @[Arbiter.scala 88:{27,36}]
  wire  _T_4 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_5 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 31:78]
  wire  _T_6 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 31:78]
  wire  _io_in_0_ready_T_1 = locked ? lockIdx == 2'h0 : 1'h1; // @[Arbiter.scala 57:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx == 2'h1 : _T_4; // @[Arbiter.scala 57:22]
  wire  _io_in_2_ready_T_1 = locked ? lockIdx == 2'h2 : _T_5; // @[Arbiter.scala 57:22]
  wire  _io_in_3_ready_T_1 = locked ? lockIdx == 2'h3 : _T_6; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_2_ready = _io_in_2_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_3_ready = _io_in_3_ready_T_1 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbiter.scala 41:{16,16}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_22; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_18; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? io_in_3_bits_cmd : _GEN_14; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_10; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_6; // @[Arbiter.scala 42:{15,15}]
  assign io_chosen = locked ? lockIdx : choice; // @[Arbiter.scala 40:13 55:{19,31}]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (_T & wantsLock) begin // @[Arbiter.scala 50:39]
      lockIdx <= io_chosen; // @[Arbiter.scala 51:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [31:0] io_in_2_req_bits_addr,
  input  [3:0]  io_in_2_req_bits_cmd,
  input  [63:0] io_in_2_req_bits_wdata,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  output        io_in_3_req_ready,
  input         io_in_3_req_valid,
  input  [31:0] io_in_3_req_bits_addr,
  input  [2:0]  io_in_3_req_bits_size,
  input  [3:0]  io_in_3_req_bits_cmd,
  input  [7:0]  io_in_3_req_bits_wmask,
  input  [63:0] io_in_3_req_bits_wdata,
  input         io_in_3_resp_ready,
  output        io_in_3_resp_valid,
  output [3:0]  io_in_3_resp_bits_cmd,
  output [63:0] io_in_3_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_3_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_3_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_3_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_3_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_3_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire [1:0] inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  reg [1:0] inflightSrc; // @[Crossbar.scala 105:24]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [1:0] _GEN_8 = _T_25 | _T_26 ? 2'h2 : state; // @[Crossbar.scala 124:{80,88} 98:22]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [1:0] _GEN_13 = _T_29 ? 2'h0 : state; // @[Crossbar.scala 128:{50,58} 98:22]
  LockingArbiter_1 inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_in_3_valid(inputArb_io_in_3_valid),
    .io_in_3_bits_addr(inputArb_io_in_3_bits_addr),
    .io_in_3_bits_size(inputArb_io_in_3_bits_size),
    .io_in_3_bits_cmd(inputArb_io_in_3_bits_cmd),
    .io_in_3_bits_wmask(inputArb_io_in_3_bits_wmask),
    .io_in_3_bits_wdata(inputArb_io_in_3_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:{13,13} 113:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = 2'h1 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:{13,13} 113:26]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[Crossbar.scala 102:68]
  assign io_in_2_resp_valid = 2'h2 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:{13,13} 113:26]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[Crossbar.scala 102:68]
  assign io_in_3_resp_valid = 2'h3 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:{13,13} 113:26]
  assign io_in_3_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[Crossbar.scala 109:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = 2'h3 == inflightSrc ? io_in_3_resp_ready : 1'h1; // @[Crossbar.scala 116:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_valid = io_in_3_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_size = io_in_3_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_cmd = io_in_3_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:37]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 98:22]
      state <= 2'h0; // @[Crossbar.scala 98:22]
    end else if (2'h0 == state) begin // @[Crossbar.scala 119:18]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        if (_T_4) begin // @[Crossbar.scala 123:38]
          state <= 2'h1; // @[Crossbar.scala 123:46]
        end else begin
          state <= _GEN_8;
        end
      end
    end else if (2'h1 == state) begin // @[Crossbar.scala 119:18]
      if (_T_29 & _T_30) begin // @[Crossbar.scala 127:82]
        state <= 2'h0; // @[Crossbar.scala 127:90]
      end
    end else if (2'h2 == state) begin // @[Crossbar.scala 119:18]
      state <= _GEN_13;
    end
    if (2'h0 == state) begin // @[Crossbar.scala 119:18]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        inflightSrc <= inputArb_io_chosen; // @[Crossbar.scala 122:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [86:0]  io_in_bits_user,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [86:0]  io_out_bits_user,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input          io_flush,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output         io_ipf,
  output         io_isFinish
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 196:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 196:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 196:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 198:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 198:30]
  wire [17:0] hi = {vpn_vpn2,vpn_vpn1}; // @[EmbeddedTLB.scala 207:201]
  wire [26:0] _T_43 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 207:201]
  wire [26:0] _T_44 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_45 = _T_44 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_47 = _T_44 & _T_43; // @[TLB.scala 131:84]
  wire  _T_48 = _T_45 == _T_47; // @[TLB.scala 131:48]
  wire  _T_49 = io_md_0[52] & io_md_0[93:78] == satp_asid & _T_48; // @[EmbeddedTLB.scala 207:132]
  wire [26:0] _T_85 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_86 = _T_85 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_88 = _T_85 & _T_43; // @[TLB.scala 131:84]
  wire  _T_89 = _T_86 == _T_88; // @[TLB.scala 131:48]
  wire  _T_90 = io_md_1[52] & io_md_1[93:78] == satp_asid & _T_89; // @[EmbeddedTLB.scala 207:132]
  wire [26:0] _T_126 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_127 = _T_126 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_129 = _T_126 & _T_43; // @[TLB.scala 131:84]
  wire  _T_130 = _T_127 == _T_129; // @[TLB.scala 131:48]
  wire  _T_131 = io_md_2[52] & io_md_2[93:78] == satp_asid & _T_130; // @[EmbeddedTLB.scala 207:132]
  wire [26:0] _T_167 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_168 = _T_167 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_170 = _T_167 & _T_43; // @[TLB.scala 131:84]
  wire  _T_171 = _T_168 == _T_170; // @[TLB.scala 131:48]
  wire  _T_172 = io_md_3[52] & io_md_3[93:78] == satp_asid & _T_171; // @[EmbeddedTLB.scala 207:132]
  wire [3:0] hitVec = {_T_172,_T_131,_T_90,_T_49}; // @[EmbeddedTLB.scala 207:211]
  wire  _T_173 = |hitVec; // @[EmbeddedTLB.scala 208:35]
  wire  hit = io_in_valid & |hitVec; // @[EmbeddedTLB.scala 208:25]
  wire  miss = io_in_valid & ~_T_173; // @[EmbeddedTLB.scala 209:26]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_182 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_185 = {_T_182,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[EmbeddedTLB.scala 211:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 212:20]
  wire [120:0] _T_192 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_193 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_194 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_195 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_196 = _T_192 | _T_193; // @[Mux.scala 27:72]
  wire [120:0] _T_197 = _T_196 | _T_194; // @[Mux.scala 27:72]
  wire [120:0] _T_198 = _T_197 | _T_195; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_198[59:52]; // @[EmbeddedTLB.scala 218:70]
  wire [17:0] hitMeta_mask = _T_198[77:60]; // @[EmbeddedTLB.scala 218:70]
  wire [15:0] hitMeta_asid = _T_198[93:78]; // @[EmbeddedTLB.scala 218:70]
  wire [31:0] hitData_pteaddr = _T_198[31:0]; // @[EmbeddedTLB.scala 219:70]
  wire [19:0] hitData_ppn = _T_198[51:32]; // @[EmbeddedTLB.scala 219:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 220:38]
  wire  _T_244 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 229:62]
  wire  _T_249 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 229:110]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u); // @[EmbeddedTLB.scala 229:87]
  wire  hitExec = hitCheck & hitFlag_x; // @[EmbeddedTLB.scala 230:26]
  wire  hitinstrPF = ~hitExec & hit; // @[EmbeddedTLB.scala 242:52]
  wire  _T_237 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 136:23]
  wire  _T_239 = ~_T_237; // @[EmbeddedTLB.scala 224:84]
  wire  hitWB = hit & ~hitFlag_a & ~hitinstrPF & ~_T_237; // @[EmbeddedTLB.scala 224:81]
  wire [7:0] _T_242 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 225:79]
  wire [7:0] hitRefillFlag = 8'h40 | _T_242; // @[EmbeddedTLB.scala 225:69]
  wire [39:0] _T_243 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 30:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  reg [2:0] state; // @[EmbeddedTLB.scala 250:22]
  reg [1:0] level; // @[EmbeddedTLB.scala 251:22]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 253:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 255:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 258:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 258:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 259:18]
  wire  _T_270 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_270 | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  reg  needFlush; // @[EmbeddedTLB.scala 263:26]
  wire  isFlush = needFlush | io_flush; // @[EmbeddedTLB.scala 265:27]
  wire  _GEN_3 = io_flush & state != 3'h0 | needFlush; // @[EmbeddedTLB.scala 263:26 266:{40,52}]
  wire  _GEN_4 = _T_270 & needFlush ? 1'h0 : _GEN_3; // @[EmbeddedTLB.scala 267:{37,49}]
  reg  missIPF; // @[EmbeddedTLB.scala 269:24]
  wire  _T_276 = ~io_flush; // @[EmbeddedTLB.scala 274:13]
  wire [31:0] _T_281 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 30:58]
  wire  _T_283 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_283 ? 3'h2 : state; // @[EmbeddedTLB.scala 250:22 291:{38,46}]
  wire  _GEN_17 = isFlush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 288:22 290:19]
  wire [7:0] _T_285 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,
    memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 295:44]
  wire  _T_294 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_297 = level == 2'h3; // @[EmbeddedTLB.scala 300:58]
  wire  _T_298 = level == 2'h2; // @[EmbeddedTLB.scala 300:73]
  wire [8:0] _T_328 = _T_297 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 314:50]
  wire [31:0] _T_330 = {memRdata_ppn,_T_328,3'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_18 = ~_T_285[0] | ~_T_285[1] & _T_285[2] ? 3'h4 : 3'h1; // @[EmbeddedTLB.scala 301:60 302:43 313:19]
  wire  _GEN_19 = ~_T_285[0] | ~_T_285[1] & _T_285[2] | missIPF; // @[EmbeddedTLB.scala 269:24 301:60 303:45]
  wire [31:0] _GEN_20 = ~_T_285[0] | ~_T_285[1] & _T_285[2] ? raddr : _T_330; // @[EmbeddedTLB.scala 259:18 301:60 314:19]
  wire  _T_343 = _T_285[0] & ~(_T_244 & ~_T_285[4]) & ~(_T_249 & _T_285[4]); // @[EmbeddedTLB.scala 317:87]
  wire  _T_344 = _T_343 & _T_285[3]; // @[EmbeddedTLB.scala 318:36]
  wire  _T_349 = ~_T_285[6]; // @[EmbeddedTLB.scala 321:60]
  wire [7:0] _T_358 = {_T_285[7],_T_285[6],_T_285[5],_T_285[4],_T_285[3],_T_285[2],_T_285[1],_T_285[0]}; // @[EmbeddedTLB.scala 323:79]
  wire [7:0] _T_359 = 8'h40 | _T_358; // @[EmbeddedTLB.scala 323:68]
  wire [63:0] _T_360 = io_mem_resp_bits_rdata | 64'h40; // @[EmbeddedTLB.scala 324:50]
  wire [2:0] _T_362 = _T_349 ? 3'h3 : 3'h4; // @[EmbeddedTLB.scala 328:27]
  wire  _GEN_21 = ~_T_344 | missIPF; // @[EmbeddedTLB.scala 269:24 326:{30,40}]
  wire [2:0] _GEN_22 = ~_T_344 ? 3'h4 : _T_362; // @[EmbeddedTLB.scala 326:{30,58} 328:21]
  wire  _GEN_23 = ~_T_344 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 326:30 329:30]
  wire [17:0] _T_365 = _T_298 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 342:59]
  wire [17:0] _T_366 = _T_297 ? 18'h0 : _T_365; // @[EmbeddedTLB.scala 342:26]
  wire [7:0] _GEN_24 = level != 2'h0 ? _T_359 : 8'h0; // @[EmbeddedTLB.scala 316:36 323:26]
  wire [63:0] _GEN_25 = level != 2'h0 ? _T_360 : memRespStore; // @[EmbeddedTLB.scala 316:36 324:24 253:25]
  wire  _GEN_26 = level != 2'h0 ? _GEN_21 : missIPF; // @[EmbeddedTLB.scala 269:24 316:36]
  wire [2:0] _GEN_27 = level != 2'h0 ? _GEN_22 : state; // @[EmbeddedTLB.scala 250:22 316:36]
  wire  _GEN_28 = level != 2'h0 & _GEN_23; // @[EmbeddedTLB.scala 316:36]
  wire [17:0] _GEN_29 = level != 2'h0 ? _T_366 : 18'h3ffff; // @[EmbeddedTLB.scala 316:36 342:20]
  wire [17:0] _GEN_37 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_29; // @[EmbeddedTLB.scala 300:82]
  wire [17:0] _GEN_45 = isFlush ? 18'h3ffff : _GEN_37; // @[EmbeddedTLB.scala 297:24]
  wire [17:0] _GEN_54 = _T_294 ? _GEN_45 : 18'h3ffff; // @[EmbeddedTLB.scala 296:33]
  wire [17:0] _GEN_77 = 3'h2 == state ? _GEN_54 : 18'h3ffff; // @[EmbeddedTLB.scala 272:18]
  wire [17:0] _GEN_88 = 3'h1 == state ? 18'h3ffff : _GEN_77; // @[EmbeddedTLB.scala 272:18]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_88; // @[EmbeddedTLB.scala 272:18]
  wire [17:0] _GEN_30 = level != 2'h0 ? missMask : missMaskStore; // @[EmbeddedTLB.scala 316:36 343:25 255:26]
  wire [2:0] _GEN_31 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_18 : _GEN_27; // @[EmbeddedTLB.scala 300:82]
  wire  _GEN_32 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_26; // @[EmbeddedTLB.scala 300:82]
  wire [31:0] _GEN_33 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : raddr; // @[EmbeddedTLB.scala 259:18 300:82]
  wire [7:0] _GEN_34 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_24; // @[EmbeddedTLB.scala 300:82]
  wire [63:0] _GEN_35 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_25; // @[EmbeddedTLB.scala 253:25 300:82]
  wire  _GEN_36 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_28; // @[EmbeddedTLB.scala 300:82]
  wire [17:0] _GEN_38 = ~(_T_285[1] | _T_285[3]) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_30; // @[EmbeddedTLB.scala 255:26 300:82]
  wire [2:0] _GEN_39 = isFlush ? 3'h0 : _GEN_31; // @[EmbeddedTLB.scala 297:24 298:17]
  wire  _GEN_40 = isFlush ? missIPF : _GEN_32; // @[EmbeddedTLB.scala 269:24 297:24]
  wire [31:0] _GEN_41 = isFlush ? raddr : _GEN_33; // @[EmbeddedTLB.scala 259:18 297:24]
  wire [7:0] _GEN_42 = isFlush ? 8'h0 : _GEN_34; // @[EmbeddedTLB.scala 297:24]
  wire [63:0] _GEN_43 = isFlush ? memRespStore : _GEN_35; // @[EmbeddedTLB.scala 297:24 253:25]
  wire  _GEN_44 = isFlush ? 1'h0 : _GEN_36; // @[EmbeddedTLB.scala 297:24]
  wire [17:0] _GEN_46 = isFlush ? missMaskStore : _GEN_38; // @[EmbeddedTLB.scala 297:24 255:26]
  wire [1:0] _T_368 = level - 2'h1; // @[EmbeddedTLB.scala 345:24]
  wire [2:0] _GEN_47 = _T_294 ? _GEN_39 : state; // @[EmbeddedTLB.scala 250:22 296:33]
  wire  _GEN_48 = _T_294 ? _GEN_17 : _GEN_4; // @[EmbeddedTLB.scala 296:33]
  wire  _GEN_49 = _T_294 ? _GEN_40 : missIPF; // @[EmbeddedTLB.scala 269:24 296:33]
  wire [7:0] _GEN_51 = _T_294 ? _GEN_42 : 8'h0; // @[EmbeddedTLB.scala 296:33]
  wire  _GEN_53 = _T_294 & _GEN_44; // @[EmbeddedTLB.scala 296:33]
  wire [1:0] _GEN_56 = _T_294 ? _T_368 : level; // @[EmbeddedTLB.scala 296:33 345:15 251:22]
  wire [2:0] _GEN_57 = _T_283 ? 3'h4 : state; // @[EmbeddedTLB.scala 250:22 353:{38,46}]
  wire [2:0] _GEN_58 = isFlush ? 3'h0 : _GEN_57; // @[EmbeddedTLB.scala 350:22 351:15]
  wire [2:0] _GEN_59 = _T_270 | io_flush | alreadyOutFire ? 3'h0 : state; // @[EmbeddedTLB.scala 356:73 357:13 250:22]
  wire  _GEN_60 = _T_270 | io_flush | alreadyOutFire ? 1'h0 : missIPF; // @[EmbeddedTLB.scala 356:73 358:15 269:24]
  wire  _GEN_61 = _T_270 | io_flush | alreadyOutFire ? 1'h0 : _GEN_2; // @[EmbeddedTLB.scala 356:73 359:22]
  wire [2:0] _GEN_62 = 3'h5 == state ? 3'h0 : state; // @[EmbeddedTLB.scala 272:18 363:13 250:22]
  wire [2:0] _GEN_63 = 3'h4 == state ? _GEN_59 : _GEN_62; // @[EmbeddedTLB.scala 272:18]
  wire  _GEN_64 = 3'h4 == state ? _GEN_60 : missIPF; // @[EmbeddedTLB.scala 272:18 269:24]
  wire  _GEN_65 = 3'h4 == state ? _GEN_61 : _GEN_2; // @[EmbeddedTLB.scala 272:18]
  wire [2:0] _GEN_66 = 3'h3 == state ? _GEN_58 : _GEN_63; // @[EmbeddedTLB.scala 272:18]
  wire  _GEN_67 = 3'h3 == state ? _GEN_17 : _GEN_4; // @[EmbeddedTLB.scala 272:18]
  wire  _GEN_68 = 3'h3 == state ? missIPF : _GEN_64; // @[EmbeddedTLB.scala 272:18 269:24]
  wire  _GEN_69 = 3'h3 == state ? _GEN_2 : _GEN_65; // @[EmbeddedTLB.scala 272:18]
  wire  _GEN_87 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_53; // @[EmbeddedTLB.scala 272:18]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_87; // @[EmbeddedTLB.scala 272:18]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 368:23]
  wire  _T_382 = ~isFlush; // @[EmbeddedTLB.scala 370:77]
  wire  _T_386 = state == 3'h0; // @[EmbeddedTLB.scala 374:82]
  reg  REG_7; // @[EmbeddedTLB.scala 374:33]
  reg [3:0] REG_9; // @[EmbeddedTLB.scala 375:60]
  reg [26:0] REG_10; // @[EmbeddedTLB.scala 375:84]
  reg [15:0] REG_11; // @[EmbeddedTLB.scala 376:19]
  reg [17:0] REG_12; // @[EmbeddedTLB.scala 376:72]
  reg [7:0] REG_13; // @[EmbeddedTLB.scala 377:19]
  reg [19:0] REG_14; // @[EmbeddedTLB.scala 377:77]
  reg [31:0] REG_15; // @[EmbeddedTLB.scala 378:22]
  wire [59:0] lo_6 = {REG_13,REG_14,REG_15}; // @[Cat.scala 30:58]
  wire [60:0] hi_13 = {REG_10,REG_11,REG_12}; // @[Cat.scala 30:58]
  wire [31:0] _T_402 = {hitData_ppn,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_404 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_405 = _T_402 & _T_404; // @[BitUtils.scala 32:13]
  wire [31:0] _T_406 = ~_T_404; // @[BitUtils.scala 32:38]
  wire [31:0] _T_407 = io_in_bits_addr[31:0] & _T_406; // @[BitUtils.scala 32:36]
  wire [31:0] _T_408 = _T_405 | _T_407; // @[BitUtils.scala 32:25]
  wire [31:0] _T_421 = {memRespStore[29:10],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_423 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_424 = _T_421 & _T_423; // @[BitUtils.scala 32:13]
  wire [31:0] _T_425 = ~_T_423; // @[BitUtils.scala 32:38]
  wire [31:0] _T_426 = io_in_bits_addr[31:0] & _T_425; // @[BitUtils.scala 32:36]
  wire [31:0] _T_427 = _T_424 | _T_426; // @[BitUtils.scala 32:25]
  wire  _T_429 = ~hitWB; // @[EmbeddedTLB.scala 383:45]
  wire  _T_436 = hit & ~hitWB ? _T_239 : state == 3'h4; // @[EmbeddedTLB.scala 383:37]
  assign io_in_ready = io_out_ready & _T_386 & ~miss & _T_429 & io_mdReady & _T_239; // @[EmbeddedTLB.scala 385:86]
  assign io_out_valid = io_in_valid & _T_436; // @[EmbeddedTLB.scala 383:31]
  assign io_out_bits_addr = hit ? _T_408 : _T_427; // @[EmbeddedTLB.scala 382:26]
  assign io_out_bits_user = io_in_bits_user; // @[EmbeddedTLB.scala 381:15]
  assign io_mdWrite_wen = REG_7; // @[TLB.scala 214:14]
  assign io_mdWrite_waymask = REG_9; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {hi_13,lo_6}; // @[Cat.scala 30:58]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~isFlush; // @[EmbeddedTLB.scala 370:74]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 369:35]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[EmbeddedTLB.scala 369:138]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 371:21]
  assign io_pf_loadPF = 1'h0; // @[EmbeddedTLB.scala 239:16]
  assign io_pf_storePF = 1'h0; // @[EmbeddedTLB.scala 240:17]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[EmbeddedTLB.scala 387:16]
  assign io_isFinish = _T_270 | _T_237; // @[EmbeddedTLB.scala 388:32]
  always @(posedge clock) begin
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_185;
    end
    if (hitWB) begin // @[Reg.scala 16:19]
      hitWBStore <= _T_243; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 250:22]
      state <= 3'h0; // @[EmbeddedTLB.scala 250:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (~io_flush & hitWB) begin // @[EmbeddedTLB.scala 274:32]
        state <= 3'h3; // @[EmbeddedTLB.scala 275:15]
      end else if (miss & _T_276) begin // @[EmbeddedTLB.scala 278:37]
        state <= 3'h1; // @[EmbeddedTLB.scala 279:15]
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (isFlush) begin // @[EmbeddedTLB.scala 288:22]
        state <= 3'h0; // @[EmbeddedTLB.scala 289:15]
      end else begin
        state <= _GEN_15;
      end
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      state <= _GEN_47;
    end else begin
      state <= _GEN_66;
    end
    if (reset) begin // @[EmbeddedTLB.scala 251:22]
      level <= 2'h3; // @[EmbeddedTLB.scala 251:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (!(~io_flush & hitWB)) begin // @[EmbeddedTLB.scala 274:32]
        if (miss & _T_276) begin // @[EmbeddedTLB.scala 278:37]
          level <= 2'h3; // @[EmbeddedTLB.scala 281:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
        level <= _GEN_56;
      end
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
          if (_T_294) begin // @[EmbeddedTLB.scala 296:33]
            memRespStore <= _GEN_43;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
          if (_T_294) begin // @[EmbeddedTLB.scala 296:33]
            missMaskStore <= _GEN_46;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (!(~io_flush & hitWB)) begin // @[EmbeddedTLB.scala 274:32]
        if (miss & _T_276) begin // @[EmbeddedTLB.scala 278:37]
          raddr <= _T_281; // @[EmbeddedTLB.scala 280:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
        if (_T_294) begin // @[EmbeddedTLB.scala 296:33]
          raddr <= _GEN_41;
        end
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (~io_flush & hitWB) begin // @[EmbeddedTLB.scala 274:32]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 277:24]
      end else if (miss & _T_276) begin // @[EmbeddedTLB.scala 278:37]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 283:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_69;
    end
    if (reset) begin // @[EmbeddedTLB.scala 263:26]
      needFlush <= 1'h0; // @[EmbeddedTLB.scala 263:26]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (~io_flush & hitWB) begin // @[EmbeddedTLB.scala 274:32]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 276:19]
      end else if (miss & _T_276) begin // @[EmbeddedTLB.scala 278:37]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 282:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (isFlush) begin // @[EmbeddedTLB.scala 288:22]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 290:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      needFlush <= _GEN_48;
    end else begin
      needFlush <= _GEN_67;
    end
    if (reset) begin // @[EmbeddedTLB.scala 269:24]
      missIPF <= 1'h0; // @[EmbeddedTLB.scala 269:24]
    end else if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
          missIPF <= _GEN_49;
        end else begin
          missIPF <= _GEN_68;
        end
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 374:33]
      REG_7 <= 1'h0; // @[EmbeddedTLB.scala 374:33]
    end else begin
      REG_7 <= missMetaRefill & _T_382 | hitWB & state == 3'h0 & _T_382; // @[EmbeddedTLB.scala 374:33]
    end
    if (hit) begin // @[EmbeddedTLB.scala 212:20]
      REG_9 <= hitVec;
    end else begin
      REG_9 <= victimWaymask;
    end
    REG_10 <= {hi,vpn_vpn0}; // @[EmbeddedTLB.scala 375:89]
    if (hitWB) begin // @[EmbeddedTLB.scala 376:23]
      REG_11 <= hitMeta_asid;
    end else begin
      REG_11 <= satp_asid;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 376:76]
      REG_12 <= hitMeta_mask;
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_12 <= 18'h3ffff;
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_12 <= 18'h3ffff;
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_12 <= _GEN_54;
    end else begin
      REG_12 <= 18'h3ffff;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 377:23]
      REG_13 <= hitRefillFlag;
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_13 <= 8'h0;
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_13 <= 8'h0;
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_13 <= _GEN_51;
    end else begin
      REG_13 <= 8'h0;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 377:81]
      REG_14 <= hitData_ppn;
    end else begin
      REG_14 <= memRdata_ppn;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 378:27]
      REG_15 <= hitData_pteaddr;
    end else begin
      REG_15 <= raddr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  hitWBStore = _RAND_1[39:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  level = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  memRespStore = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  missMaskStore = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  raddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  alreadyOutFire = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  needFlush = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  missIPF = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_9 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  REG_10 = _RAND_12[26:0];
  _RAND_13 = {1{`RANDOM}};
  REG_11 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  REG_12 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  REG_13 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  REG_14 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  REG_15 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_1 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_2 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_3 [0:0]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg  resetState; // @[EmbeddedTLB.scala 55:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[EmbeddedTLB.scala 57:22 55:27 57:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 66:20]
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = 1'h0;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = 1'h0;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = 1'h0;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = 1'h0;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = 1'h0;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = 1'h0;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = 1'h0;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = 1'h0;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 72:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    resetState <= reset | _GEN_1; // @[EmbeddedTLB.scala 55:{27,27}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [86:0] io_out_req_bits_user,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input  [86:0] io_out_resp_bits_user,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_flush,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_cacheEmpty,
  output        io_ipf,
  input  [63:0] CSRSATP,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 83:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 83:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 83:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 83:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 83:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 83:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 83:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_flush; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 83:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_ipf; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 83:23]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 85:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 85:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 85:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 85:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 85:21]
  reg [120:0] r__0; // @[Reg.scala 15:16]
  reg [120:0] r__1; // @[Reg.scala 15:16]
  reg [120:0] r__2; // @[Reg.scala 15:16]
  reg [120:0] r__3; // @[Reg.scala 15:16]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 117:26]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 105:57]
  reg  REG; // @[EmbeddedTLB.scala 108:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : REG; // @[EmbeddedTLB.scala 108:24 109:{25,33}]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[EmbeddedTLB.scala 110:{50,58}]
  reg [38:0] r_1_addr; // @[Reg.scala 15:16]
  reg [86:0] r_1_user; // @[Reg.scala 15:16]
  wire  _GEN_13 = ~vmEnable | io_out_req_ready; // @[EmbeddedTLB.scala 126:19 127:26 139:23]
  wire  _GEN_14 = ~vmEnable ? io_in_req_valid : tlbExec_io_out_valid; // @[EmbeddedTLB.scala 126:19 129:22 139:23]
  wire  _T_17 = tlbExec_io_ipf & vmEnable; // @[EmbeddedTLB.scala 155:26]
  EmbeddedTLBExec tlbExec ( // @[EmbeddedTLB.scala 83:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish)
  );
  EmbeddedTLBMD mdTLB ( // @[EmbeddedTLB.scala 85:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 113:16 126:19 130:21]
  assign io_in_resp_valid = _T_17 & io_cacheEmpty | io_out_resp_valid; // @[EmbeddedTLB.scala 141:15 160:56 161:24]
  assign io_in_resp_bits_rdata = _T_17 & io_cacheEmpty ? 64'h0 : io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 141:15 160:56 162:29]
  assign io_in_resp_bits_user = _T_17 & io_cacheEmpty ? tlbExec_io_in_bits_user : io_out_resp_bits_user; // @[EmbeddedTLB.scala 141:15 160:56 164:34]
  assign io_out_req_valid = tlbExec_io_ipf & vmEnable ? 1'h0 : _GEN_14; // @[EmbeddedTLB.scala 155:39 157:24]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 126:19 131:26 139:23]
  assign io_out_req_bits_user = ~vmEnable ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 126:19 136:32 139:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[EmbeddedTLB.scala 141:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 90:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 90:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 90:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 90:18]
  assign io_ipf = _T_17 & io_cacheEmpty & tlbExec_io_ipf; // @[EmbeddedTLB.scala 160:56 165:14 97:10]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = REG; // @[EmbeddedTLB.scala 115:17]
  assign tlbExec_io_in_bits_addr = r_1_addr; // @[EmbeddedTLB.scala 114:16]
  assign tlbExec_io_in_bits_user = r_1_user; // @[EmbeddedTLB.scala 114:16]
  assign tlbExec_io_out_ready = tlbExec_io_ipf & vmEnable ? io_cacheEmpty & io_in_resp_ready : _GEN_13; // @[EmbeddedTLB.scala 155:39 156:28]
  assign tlbExec_io_md_0 = r__0; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_md_1 = r__1; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_md_2 = r__2; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_md_3 = r__3; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 93:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 90:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 90:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 90:18]
  assign tlbExec_io_flush = io_flush; // @[EmbeddedTLB.scala 88:20]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 89:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 91:17]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 102:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 95:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 95:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 95:18]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__0 <= mdTLB_io_tlbmd_0; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__1 <= mdTLB_io_tlbmd_1; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__2 <= mdTLB_io_tlbmd_2; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__3 <= mdTLB_io_tlbmd_3; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 108:24]
      REG <= 1'h0; // @[EmbeddedTLB.scala 108:24]
    end else if (io_flush) begin // @[EmbeddedTLB.scala 111:20]
      REG <= 1'h0; // @[EmbeddedTLB.scala 111:28]
    end else begin
      REG <= _GEN_5;
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r_1_addr <= io_in_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r_1_user <= io_in_req_bits_user; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  r__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  r__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  r__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  r__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  r_1_addr = _RAND_5[38:0];
  _RAND_6 = {3{`RANDOM}};
  r_1_user = _RAND_6[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [86:0] io_in_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [86:0] io_out_bits_req_user,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_22 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_22) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 147:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 146:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 145:19]
  assign io_out_bits_req_user = io_in_bits_user; // @[Cache.scala 145:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module CacheStage2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [86:0] io_in_bits_req_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [86:0] io_out_bits_req_user,
  output [18:0] io_out_bits_metas_0_tag,
  output [18:0] io_out_bits_metas_1_tag,
  output [18:0] io_out_bits_metas_2_tag,
  output [18:0] io_out_bits_metas_3_tag,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 176:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 176:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 176:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 178:64]
  reg  isForwardMetaReg; // @[Cache.scala 179:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 180:24 179:33 180:43]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 181:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 181:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 15:16 16:{19,23}]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 15:16 16:{19,23}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 185:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 187:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 187:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 187:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 187:61]
  wire [18:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[Cache.scala 189:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 192:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_39 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_42 = {_T_39,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 193:42]
  wire  _T_45 = ~metaWay_0_valid; // @[Cache.scala 195:45]
  wire  _T_46 = ~metaWay_1_valid; // @[Cache.scala 195:45]
  wire  _T_47 = ~metaWay_2_valid; // @[Cache.scala 195:45]
  wire  _T_48 = ~metaWay_3_valid; // @[Cache.scala 195:45]
  wire [3:0] invalidVec = {_T_48,_T_47,_T_46,_T_45}; // @[Cache.scala 195:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 196:34]
  wire [1:0] _T_52 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 199:8]
  wire [2:0] _T_53 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_52}; // @[Cache.scala 198:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_53}; // @[Cache.scala 197:33]
  wire [3:0] _T_54 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 202:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  wire [1:0] _T_59 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_61 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_63 = _T_59 + _T_61; // @[Bitwise.scala 47:55]
  wire  _T_65 = _T_63 > 3'h1; // @[Cache.scala 203:26]
  wire [31:0] _T_172 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 87:11]
  wire  _T_174 = _T_172[31:28] == 4'h0; // @[NutCore.scala 87:44]
  wire [31:0] _T_175 = io_in_bits_req_addr ^ 32'h40600000; // @[NutCore.scala 87:11]
  wire  _T_177 = _T_175[31:24] == 8'h0; // @[NutCore.scala 87:44]
  wire [9:0] _T_187 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_189 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_187; // @[Cache.scala 219:13]
  wire  isForwardData = io_in_valid & _T_189; // @[Cache.scala 218:35]
  reg  isForwardDataReg; // @[Cache.scala 221:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 222:24 221:33 222:43]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_196 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_196; // @[Cache.scala 230:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 229:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 228:19]
  assign io_out_bits_req_user = io_in_bits_req_user; // @[Cache.scala 228:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 215:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 213:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  assign io_out_bits_mmio = _T_174 | _T_177; // @[NutCore.scala 88:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 225:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 226:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 226:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 179:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 179:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 181:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 181:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_42;
    end
    if (reset) begin // @[Cache.scala 221:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 221:33]
    end else if (_T_12) begin // @[Cache.scala 223:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 223:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 16:23]
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:210 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 210:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fatal; // @[Cache.scala 210:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  REG = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  isForwardDataReg = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_6[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  input         io_in_0_valid,
  input  [6:0]  io_in_0_bits_setIdx,
  input  [18:0] io_in_0_bits_data_tag,
  input         io_in_0_bits_data_dirty,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [6:0]  io_in_1_bits_setIdx,
  input  [18:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [6:0]  io_out_bits_setIdx,
  output [18:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid ? io_in_0_bits_data_dirty : io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module Arbiter_1(
  input         io_in_0_valid,
  input  [9:0]  io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [9:0]  io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [9:0]  io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module CacheStage3(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [86:0] io_in_bits_req_user,
  input  [18:0] io_in_bits_metas_0_tag,
  input  [18:0] io_in_bits_metas_1_tag,
  input  [18:0] io_in_bits_metas_2_tag,
  input  [18:0] io_in_bits_metas_3_tag,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_rdata,
  output [86:0] io_out_bits_user,
  output        io_isFinish,
  input         io_flush,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 256:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 256:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 256:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 256:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 256:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 256:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 256:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 257:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 257:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 257:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 257:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 260:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 260:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 261:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 262:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 263:26]
  wire [18:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [18:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 275:49]
  wire [63:0] _T_43 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_43 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_48 | _T_46; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_49; // @[Cache.scala 277:21]
  wire  _T_78 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [3:0] state; // @[Cache.scala 296:22]
  reg  needFlush; // @[Cache.scala 297:26]
  wire  _GEN_1 = io_flush & state != 4'h0 | needFlush; // @[Cache.scala 297:26 299:{41,53}]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 306:23]
  wire  _T_103 = state == 4'h3; // @[Cache.scala 308:39]
  wire  _T_104 = state == 4'h8; // @[Cache.scala 308:66]
  wire [2:0] _T_109 = _T_104 ? value_1 : value_2; // @[Cache.scala 309:33]
  wire  _T_111 = state2 == 2'h1; // @[Cache.scala 310:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_116 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_117 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_118 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_119 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_120 = _T_116 | _T_117; // @[Mux.scala 27:72]
  wire [63:0] _T_121 = _T_120 | _T_118; // @[Mux.scala 27:72]
  wire  _T_124 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_127 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_8 = _T_127 | io_cohResp_valid ? 2'h0 : state2; // @[Cache.scala 316:{100,109} 306:23]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_133 = state == 4'h1; // @[Cache.scala 324:23]
  wire [2:0] _T_135 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 325:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_135; // @[Cache.scala 324:16]
  wire  _T_141 = state2 == 2'h2; // @[Cache.scala 331:89]
  reg  afterFirstRead; // @[Cache.scala 338:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_78 | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  wire  _T_147 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_149 = state == 4'h2; // @[Cache.scala 340:70]
  wire  readingFirst = ~afterFirstRead & _T_147 & state == 4'h2; // @[Cache.scala 340:60]
  wire  _T_152 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 342:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_153 = state == 4'h0; // @[Cache.scala 345:31]
  wire  _T_187 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_189 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = _T_189 ? 4'h7 : state; // @[Cache.scala 296:22 374:{50,58}]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid ? _value_T_7 : value_1; // @[Cache.scala 377:48 Counter.scala 76:15 60:40]
  wire [3:0] _GEN_29 = _T_127 ? 4'h2 : state; // @[Cache.scala 381:50 382:13 296:22]
  wire [2:0] _GEN_30 = _T_127 ? addr_wordIndex : value_1; // @[Cache.scala 381:50 383:25 Counter.scala 60:40]
  wire  _T_203 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_203 ? 4'h7 : state; // @[Cache.scala 296:22 391:{46,54}]
  wire  _GEN_33 = _T_147 | afterFirstRead; // @[Cache.scala 387:33 388:24 338:31]
  wire [2:0] _GEN_34 = _T_147 ? _value_T_7 : value_1; // @[Cache.scala 387:33 Counter.scala 76:15 60:40]
  wire [3:0] _GEN_36 = _T_147 ? _GEN_32 : state; // @[Cache.scala 296:22 387:33]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_127 ? _value_T_11 : value_2; // @[Cache.scala 396:32 Counter.scala 76:15 60:40]
  wire  _T_206 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_206 & _T_127 ? 4'h4 : state; // @[Cache.scala 296:22 397:{65,73}]
  wire [3:0] _GEN_39 = _T_147 ? 4'h1 : state; // @[Cache.scala 296:22 400:{53,61}]
  wire [3:0] _GEN_40 = _T_78 | needFlush | alreadyOutFire ? 4'h0 : state; // @[Cache.scala 296:22 401:{76,84}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[Cache.scala 355:18 296:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[Cache.scala 355:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : value_2; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[Cache.scala 355:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : value_1; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[Cache.scala 355:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? value_2 : _GEN_43; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[Cache.scala 355:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[Cache.scala 355:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_54 = 4'h1 == state ? value_2 : _GEN_49; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[Cache.scala 355:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? state : _GEN_50; // @[Cache.scala 355:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_59 = 4'h8 == state ? value_2 : _GEN_54; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire  dataRefillWriteBus_req_valid = _T_149 & _T_147; // @[Cache.scala 406:39]
  wire  _T_248 = state == 4'h7; // @[Cache.scala 448:48]
  wire  _T_267 = mmio ? _T_248 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 449:45]
  wire  _T_268 = hit | _T_267; // @[Cache.scala 449:28]
  Arbiter metaWriteArb ( // @[Cache.scala 256:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 257:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & _T_153 & ~miss; // @[Cache.scala 460:70]
  assign io_out_valid = io_in_valid & _T_268; // @[Cache.scala 447:31]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 441:29]
  assign io_out_bits_user = io_in_bits_req_user; // @[Cache.scala 444:56]
  assign io_isFinish = hit ? _T_78 : _T_248 & _GEN_12; // @[Cache.scala 457:8]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 308:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_109}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 411:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 421:23]
  assign io_mem_req_valid = _T_133 | _T_103 & state2 == 2'h2; // @[Cache.scala 331:48]
  assign io_mem_req_bits_addr = _T_133 ? raddr : waddr; // @[Cache.scala 326:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_121 | _T_119; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 330:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 336:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 334:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 335:22]
  assign io_cohResp_valid = _T_104 & _T_141; // @[Cache.scala 346:46]
  assign metaWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 291:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h0; // @[Cache.scala 292:16 97:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 290:29 SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_203; // @[Cache.scala 414:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 260:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = 1'h0; // @[Cache.scala 415:85]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 413:32 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 285:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = useForwardData ? io_in_bits_forwardData_data_data : _T_49; // @[Cache.scala 277:21]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 286:29 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _T_149 & _T_147; // @[Cache.scala 406:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = io_mem_resp_bits_rdata; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:32 SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 296:22]
      state <= 4'h0; // @[Cache.scala 296:22]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      if ((miss | mmio) & ~io_flush) begin // @[Cache.scala 368:49]
        if (mmio) begin // @[Cache.scala 369:21]
          state <= 4'h5;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (4'h5 == state) begin // @[Cache.scala 355:18]
      if (_T_187) begin // @[Cache.scala 373:48]
        state <= 4'h6; // @[Cache.scala 373:56]
      end
    end else if (4'h6 == state) begin // @[Cache.scala 355:18]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[Cache.scala 297:26]
      needFlush <= 1'h0; // @[Cache.scala 297:26]
    end else if (_T_78 & needFlush) begin // @[Cache.scala 300:37]
      needFlush <= 1'h0; // @[Cache.scala 300:49]
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
          value_1 <= _GEN_55;
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 306:23]
      state2 <= 2'h0; // @[Cache.scala 306:23]
    end else if (2'h0 == state2) begin // @[Cache.scala 313:19]
      if (_T_124) begin // @[Cache.scala 314:53]
        state2 <= 2'h1; // @[Cache.scala 314:62]
      end
    end else if (2'h1 == state2) begin // @[Cache.scala 313:19]
      state2 <= 2'h2; // @[Cache.scala 315:35]
    end else if (2'h2 == state2) begin // @[Cache.scala 313:19]
      state2 <= _GEN_8;
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Cache.scala 338:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 338:31]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      afterFirstRead <= 1'h0; // @[Cache.scala 357:22]
    end else if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      alreadyOutFire <= 1'h0; // @[Cache.scala 358:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_152) begin // @[Reg.scala 16:19]
      if (mmio) begin // @[Cache.scala 341:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:267 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 267:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 267:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  needFlush = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_1(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [6:0]  io_rreq_bits_setIdx,
  output [18:0] io_rresp_data_0_tag,
  output        io_rresp_data_0_valid,
  output        io_rresp_data_0_dirty,
  output [18:0] io_rresp_data_1_tag,
  output        io_rresp_data_1_valid,
  output        io_rresp_data_1_dirty,
  output [18:0] io_rresp_data_2_tag,
  output        io_rresp_data_2_valid,
  output        io_rresp_data_2_dirty,
  output [18:0] io_rresp_data_3_tag,
  output        io_rresp_data_3_valid,
  output        io_rresp_data_3_dirty,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [18:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  reg  REG; // @[SRAMTemplate.scala 80:30]
  reg [6:0] value; // @[Counter.scala 60:40]
  wire  wrap_wrap = value == 7'h7f; // @[Counter.scala 72:24]
  wire [6:0] _wrap_value_T_1 = value + 7'h1; // @[Counter.scala 76:24]
  wire  wrap = REG & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = wrap ? 1'h0 : REG; // @[SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  wire  _T = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
  wire [6:0] setIdx = REG ? value : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [20:0] _T_1 = {io_wreq_bits_data_tag,1'h1,io_wreq_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = REG ? 4'hf : io_wreq_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [20:0] _WIRE_2 = array_RW0_rdata_0;
  wire [20:0] _WIRE_3 = array_RW0_rdata_1;
  wire [20:0] _WIRE_4 = array_RW0_rdata_2;
  wire [20:0] _WIRE_5 = array_RW0_rdata_3;
  array_0 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~REG & _T; // @[SRAMTemplate.scala 101:33]
  assign io_rresp_data_0_tag = _WIRE_2[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_valid = _WIRE_2[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_dirty = _WIRE_2[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_tag = _WIRE_3[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_valid = _WIRE_3[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_dirty = _WIRE_3[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_tag = _WIRE_4[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_valid = _WIRE_4[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_dirty = _WIRE_4[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_tag = _WIRE_5[20:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_valid = _WIRE_5[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_dirty = _WIRE_5[0]; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = REG ? 21'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | wen;
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[Counter.scala 60:40]
      value <= 7'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      value <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_2(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [6:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [6:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [6:0]  io_r0_req_bits_setIdx,
  output [18:0] io_r0_resp_data_0_tag,
  output        io_r0_resp_data_0_valid,
  output        io_r0_resp_data_0_dirty,
  output [18:0] io_r0_resp_data_1_tag,
  output        io_r0_resp_data_1_valid,
  output        io_r0_resp_data_1_dirty,
  output [18:0] io_r0_resp_data_2_tag,
  output        io_r0_resp_data_2_valid,
  output        io_r0_resp_data_2_dirty,
  output [18:0] io_r0_resp_data_3_tag,
  output        io_r0_resp_data_3_valid,
  output        io_r0_resp_data_3_dirty,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [18:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_wreq_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [18:0] r_0_tag; // @[Reg.scala 27:20]
  reg  r_0_valid; // @[Reg.scala 27:20]
  reg  r_0_dirty; // @[Reg.scala 27:20]
  reg [18:0] r_1_tag; // @[Reg.scala 27:20]
  reg  r_1_valid; // @[Reg.scala 27:20]
  reg  r_1_dirty; // @[Reg.scala 27:20]
  reg [18:0] r_2_tag; // @[Reg.scala 27:20]
  reg  r_2_valid; // @[Reg.scala 27:20]
  reg  r_2_dirty; // @[Reg.scala 27:20]
  reg [18:0] r_3_tag; // @[Reg.scala 27:20]
  reg  r_3_valid; // @[Reg.scala 27:20]
  reg  r_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_1 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(ram_io_rresp_data_0_tag),
    .io_rresp_data_0_valid(ram_io_rresp_data_0_valid),
    .io_rresp_data_0_dirty(ram_io_rresp_data_0_dirty),
    .io_rresp_data_1_tag(ram_io_rresp_data_1_tag),
    .io_rresp_data_1_valid(ram_io_rresp_data_1_valid),
    .io_rresp_data_1_dirty(ram_io_rresp_data_1_dirty),
    .io_rresp_data_2_tag(ram_io_rresp_data_2_tag),
    .io_rresp_data_2_valid(ram_io_rresp_data_2_valid),
    .io_rresp_data_2_dirty(ram_io_rresp_data_2_dirty),
    .io_rresp_data_3_tag(ram_io_rresp_data_3_tag),
    .io_rresp_data_3_valid(ram_io_rresp_data_3_valid),
    .io_rresp_data_3_dirty(ram_io_rresp_data_3_dirty),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(ram_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(ram_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_2 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_tag = REG ? ram_io_rresp_data_0_tag : r_0_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_valid = REG ? ram_io_rresp_data_0_valid : r_0_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_dirty = REG ? ram_io_rresp_data_0_dirty : r_0_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_tag = REG ? ram_io_rresp_data_1_tag : r_1_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_valid = REG ? ram_io_rresp_data_1_valid : r_1_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_dirty = REG ? ram_io_rresp_data_1_dirty : r_1_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_tag = REG ? ram_io_rresp_data_2_tag : r_2_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_valid = REG ? ram_io_rresp_data_2_valid : r_2_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_dirty = REG ? ram_io_rresp_data_2_dirty : r_2_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_tag = REG ? ram_io_rresp_data_3_tag : r_3_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_valid = REG ? ram_io_rresp_data_3_valid : r_3_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_dirty = REG ? ram_io_rresp_data_3_dirty : r_3_dirty; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_tag = io_wreq_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_dirty = io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_0_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_tag <= ram_io_rresp_data_0_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_valid <= ram_io_rresp_data_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_dirty <= ram_io_rresp_data_0_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_tag <= ram_io_rresp_data_1_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_valid <= ram_io_rresp_data_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_dirty <= ram_io_rresp_data_1_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_tag <= ram_io_rresp_data_2_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_valid <= ram_io_rresp_data_2_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_dirty <= ram_io_rresp_data_2_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_tag <= 19'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_tag <= ram_io_rresp_data_3_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_valid <= ram_io_rresp_data_3_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_dirty <= ram_io_rresp_data_3_dirty; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_0_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  r_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1_tag = _RAND_4[18:0];
  _RAND_5 = {1{`RANDOM}};
  r_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_2_tag = _RAND_7[18:0];
  _RAND_8 = {1{`RANDOM}};
  r_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_3_tag = _RAND_10[18:0];
  _RAND_11 = {1{`RANDOM}};
  r_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_2(
  input         clock,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [9:0]  io_rreq_bits_setIdx,
  output [63:0] io_rresp_data_0_data,
  output [63:0] io_rresp_data_1_data,
  output [63:0] io_rresp_data_2_data,
  output [63:0] io_rresp_data_3_data,
  input         io_wreq_valid,
  input  [9:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
  wire [9:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  wire  realRen = io_rreq_valid & ~io_wreq_valid; // @[SRAMTemplate.scala 89:38]
  array_1 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~io_wreq_valid; // @[SRAMTemplate.scala 101:53]
  assign io_rresp_data_0_data = array_RW0_rdata_0; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_data = array_RW0_rdata_1; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_data = array_RW0_rdata_2; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_data = array_RW0_rdata_3; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = io_wreq_bits_waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = io_wreq_bits_waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = io_wreq_bits_waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = io_wreq_bits_waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | io_wreq_valid;
  assign array_RW0_wmode = io_wreq_valid; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx;
endmodule
module Arbiter_3(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [9:0] io_in_0_bits_setIdx,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [9:0] io_in_1_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [9:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module SRAMTemplateWithArbiter_1(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [9:0]  io_r0_req_bits_setIdx,
  output [63:0] io_r0_resp_data_0_data,
  output [63:0] io_r0_resp_data_1_data,
  output [63:0] io_r0_resp_data_2_data,
  output [63:0] io_r0_resp_data_3_data,
  output        io_r1_req_ready,
  input         io_r1_req_valid,
  input  [9:0]  io_r1_req_bits_setIdx,
  output [63:0] io_r1_resp_data_0_data,
  output [63:0] io_r1_resp_data_1_data,
  output [63:0] io_r1_resp_data_2_data,
  output [63:0] io_r1_resp_data_3_data,
  input         io_wreq_valid,
  input  [9:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_wreq_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r__0_data; // @[Reg.scala 27:20]
  reg [63:0] r__1_data; // @[Reg.scala 27:20]
  reg [63:0] r__2_data; // @[Reg.scala 27:20]
  reg [63:0] r__3_data; // @[Reg.scala 27:20]
  reg  REG_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r_1_0_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_1_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_2_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_2 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_data(ram_io_rresp_data_0_data),
    .io_rresp_data_1_data(ram_io_rresp_data_1_data),
    .io_rresp_data_2_data(ram_io_rresp_data_2_data),
    .io_rresp_data_3_data(ram_io_rresp_data_3_data),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(ram_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_3 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_data = REG ? ram_io_rresp_data_0_data : r__0_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_data = REG ? ram_io_rresp_data_1_data : r__1_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_data = REG ? ram_io_rresp_data_2_data : r__2_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_data = REG ? ram_io_rresp_data_3_data : r__3_data; // @[Hold.scala 23:48]
  assign io_r1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r1_resp_data_0_data = REG_1 ? ram_io_rresp_data_0_data : r_1_0_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_1_data = REG_1 ? ram_io_rresp_data_1_data : r_1_1_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_2_data = REG_1 ? ram_io_rresp_data_2_data : r_1_2_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_3_data = REG_1 ? ram_io_rresp_data_3_data : r_1_3_data; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_data = io_wreq_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r__0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
    REG_1 <= io_r1_req_ready & io_r1_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_1_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r__0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r__1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  r__2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  r__3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r_1_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  r_1_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  r_1_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_4(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [86:0] io_in_0_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [86:0] io_out_bits_user
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[Arbiter.scala 124:15]
  assign io_out_bits_user = io_in_0_bits_user; // @[Arbiter.scala 124:15]
endmodule
module Cache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input  [1:0]  io_flush,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_empty,
  input         MOUFlushICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 482:18]
  wire  s1_io_in_valid; // @[Cache.scala 482:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 482:18]
  wire [86:0] s1_io_in_bits_user; // @[Cache.scala 482:18]
  wire  s1_io_out_ready; // @[Cache.scala 482:18]
  wire  s1_io_out_valid; // @[Cache.scala 482:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 482:18]
  wire [86:0] s1_io_out_bits_req_user; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 482:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 482:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 482:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 482:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 482:18]
  wire  s2_clock; // @[Cache.scala 483:18]
  wire  s2_reset; // @[Cache.scala 483:18]
  wire  s2_io_in_ready; // @[Cache.scala 483:18]
  wire  s2_io_in_valid; // @[Cache.scala 483:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 483:18]
  wire [86:0] s2_io_in_bits_req_user; // @[Cache.scala 483:18]
  wire  s2_io_out_ready; // @[Cache.scala 483:18]
  wire  s2_io_out_valid; // @[Cache.scala 483:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 483:18]
  wire [86:0] s2_io_out_bits_req_user; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 483:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 483:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 483:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 483:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 483:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 483:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 483:18]
  wire  s3_clock; // @[Cache.scala 484:18]
  wire  s3_reset; // @[Cache.scala 484:18]
  wire  s3_io_in_ready; // @[Cache.scala 484:18]
  wire  s3_io_in_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 484:18]
  wire [86:0] s3_io_in_bits_req_user; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 484:18]
  wire  s3_io_out_ready; // @[Cache.scala 484:18]
  wire  s3_io_out_valid; // @[Cache.scala 484:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 484:18]
  wire [86:0] s3_io_out_bits_user; // @[Cache.scala 484:18]
  wire  s3_io_isFinish; // @[Cache.scala 484:18]
  wire  s3_io_flush; // @[Cache.scala 484:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 484:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 484:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 484:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 484:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 484:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 484:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 484:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 484:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 484:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 484:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 484:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 484:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 484:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 484:18]
  wire  metaArray_clock; // @[Cache.scala 485:25]
  wire  metaArray_reset; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 485:25]
  wire [6:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 485:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 485:25]
  wire [6:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 485:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 485:25]
  wire  dataArray_clock; // @[Cache.scala 486:25]
  wire  dataArray_reset; // @[Cache.scala 486:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 486:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 486:25]
  wire [9:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 486:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 486:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 486:25]
  wire [9:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 486:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 486:25]
  wire [9:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 486:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 486:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 495:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 495:19]
  wire [86:0] arb_io_in_0_bits_user; // @[Cache.scala 495:19]
  wire  arb_io_out_ready; // @[Cache.scala 495:19]
  wire  arb_io_out_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 495:19]
  wire [86:0] arb_io_out_bits_user; // @[Cache.scala 495:19]
  wire  _T_2 = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_2 ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_4 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_req_addr; // @[Reg.scala 15:16]
  reg [86:0] r_req_user; // @[Reg.scala 15:16]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_9 = s3_io_isFinish ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_7 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_10 = s2_io_out_valid & s3_io_in_ready | _GEN_9; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [86:0] r_1_req_user; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_0_tag; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_1_tag; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_2_tag; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_3_tag; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_3_data; // @[Reg.scala 15:16]
  reg  r_1_hit; // @[Reg.scala 15:16]
  reg [3:0] r_1_waymask; // @[Reg.scala 15:16]
  reg  r_1_mmio; // @[Reg.scala 15:16]
  reg  r_1_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] r_1_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] r_1_forwardData_waymask; // @[Reg.scala 15:16]
  CacheStage1 s1 ( // @[Cache.scala 482:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_user(s1_io_in_bits_user),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_user(s1_io_out_bits_req_user),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2 s2 ( // @[Cache.scala 483:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_user(s2_io_in_bits_req_user),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_user(s2_io_out_bits_req_user),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3 s3 ( // @[Cache.scala 484:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_user(s3_io_in_bits_req_user),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_out_bits_user(s3_io_out_bits_user),
    .io_isFinish(s3_io_isFinish),
    .io_flush(s3_io_flush),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 485:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 486:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_4 arb ( // @[Cache.scala 495:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_user(arb_io_in_0_bits_user),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_user(arb_io_out_bits_user)
  );
  assign io_in_req_ready = arb_io_in_0_ready; // @[Cache.scala 496:28]
  assign io_in_resp_valid = s3_io_out_valid; // @[Cache.scala 512:100]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 506:14]
  assign io_in_resp_bits_user = s3_io_out_bits_user; // @[Cache.scala 506:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 508:14]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 509:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 509:11]
  assign io_empty = ~s2_io_in_valid & ~s3_io_in_valid; // @[Cache.scala 510:31]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 498:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 498:12]
  assign s1_io_in_bits_user = arb_io_out_bits_user; // @[Cache.scala 498:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 530:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 531:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = r_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_user = r_req_user; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 537:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 540:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 539:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = r_1_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_user = r_1_req_user; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = r_1_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = r_1_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = r_1_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = r_1_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = r_1_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = r_1_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = r_1_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = r_1_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = r_1_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = r_1_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = r_1_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = r_1_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = r_1_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = r_1_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 506:14]
  assign s3_io_flush = io_flush[1]; // @[Cache.scala 507:26]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 532:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 508:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 509:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 509:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 509:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset | MOUFlushICache; // @[Cache.scala 492:37]
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 530:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 530:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 534:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 531:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 531:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 532:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 532:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 535:18]
  assign arb_io_in_0_valid = io_in_req_valid; // @[Cache.scala 496:28]
  assign arb_io_in_0_bits_addr = io_in_req_bits_addr; // @[Cache.scala 496:28]
  assign arb_io_in_0_bits_user = io_in_req_bits_user; // @[Cache.scala 496:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 498:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_4) begin // @[Reg.scala 16:19]
      r_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_4) begin // @[Reg.scala 16:19]
      r_req_user <= s1_io_out_bits_req_user; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[Pipeline.scala 27:20]
      REG_1 <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG_1 <= _GEN_10;
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_req_user <= s2_io_out_bits_req_user; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_hit <= s2_io_out_bits_hit; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 16:23]
    end
    if (_T_7) begin // @[Reg.scala 16:19]
      r_1_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_req_addr = _RAND_1[31:0];
  _RAND_2 = {3{`RANDOM}};
  r_req_user = _RAND_2[86:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1_req_addr = _RAND_4[31:0];
  _RAND_5 = {3{`RANDOM}};
  r_1_req_user = _RAND_5[86:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_metas_0_tag = _RAND_6[18:0];
  _RAND_7 = {1{`RANDOM}};
  r_1_metas_1_tag = _RAND_7[18:0];
  _RAND_8 = {1{`RANDOM}};
  r_1_metas_2_tag = _RAND_8[18:0];
  _RAND_9 = {1{`RANDOM}};
  r_1_metas_3_tag = _RAND_9[18:0];
  _RAND_10 = {2{`RANDOM}};
  r_1_datas_0_data = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  r_1_datas_1_data = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  r_1_datas_2_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  r_1_datas_3_data = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  r_1_hit = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_1_waymask = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_mmio = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_1_isForwardData = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  r_1_forwardData_data_data = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  r_1_forwardData_waymask = _RAND_19[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [2:0]   io_in_bits_size,
  input  [3:0]   io_in_bits_cmd,
  input  [7:0]   io_in_bits_wmask,
  input  [63:0]  io_in_bits_wdata,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_cmd,
  output [7:0]   io_out_bits_wmask,
  output [63:0]  io_out_bits_wdata,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_windex,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  input          io_pf_status_sum,
  input          io_pf_status_mxr,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output [38:0]  io_pf_addr,
  output         io_isFinish,
  input          ISAMO
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 196:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 196:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 196:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 198:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 198:30]
  wire [17:0] hi = {vpn_vpn2,vpn_vpn1}; // @[EmbeddedTLB.scala 207:201]
  wire [26:0] _T_43 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 207:201]
  wire [26:0] _T_44 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_45 = _T_44 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_47 = _T_44 & _T_43; // @[TLB.scala 131:84]
  wire  _T_48 = _T_45 == _T_47; // @[TLB.scala 131:48]
  wire  _T_49 = io_md_0[52] & io_md_0[93:78] == satp_asid & _T_48; // @[EmbeddedTLB.scala 207:132]
  wire [26:0] _T_85 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_86 = _T_85 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_88 = _T_85 & _T_43; // @[TLB.scala 131:84]
  wire  _T_89 = _T_86 == _T_88; // @[TLB.scala 131:48]
  wire  _T_90 = io_md_1[52] & io_md_1[93:78] == satp_asid & _T_89; // @[EmbeddedTLB.scala 207:132]
  wire [26:0] _T_126 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_127 = _T_126 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_129 = _T_126 & _T_43; // @[TLB.scala 131:84]
  wire  _T_130 = _T_127 == _T_129; // @[TLB.scala 131:48]
  wire  _T_131 = io_md_2[52] & io_md_2[93:78] == satp_asid & _T_130; // @[EmbeddedTLB.scala 207:132]
  wire [26:0] _T_167 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_168 = _T_167 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_170 = _T_167 & _T_43; // @[TLB.scala 131:84]
  wire  _T_171 = _T_168 == _T_170; // @[TLB.scala 131:48]
  wire  _T_172 = io_md_3[52] & io_md_3[93:78] == satp_asid & _T_171; // @[EmbeddedTLB.scala 207:132]
  wire [3:0] hitVec = {_T_172,_T_131,_T_90,_T_49}; // @[EmbeddedTLB.scala 207:211]
  wire  _T_173 = |hitVec; // @[EmbeddedTLB.scala 208:35]
  wire  hit = io_in_valid & |hitVec; // @[EmbeddedTLB.scala 208:25]
  wire  miss = io_in_valid & ~_T_173; // @[EmbeddedTLB.scala 209:26]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_182 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_185 = {_T_182,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[EmbeddedTLB.scala 211:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 212:20]
  wire [120:0] _T_192 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_193 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_194 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_195 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_196 = _T_192 | _T_193; // @[Mux.scala 27:72]
  wire [120:0] _T_197 = _T_196 | _T_194; // @[Mux.scala 27:72]
  wire [120:0] _T_198 = _T_197 | _T_195; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_198[59:52]; // @[EmbeddedTLB.scala 218:70]
  wire [17:0] hitMeta_mask = _T_198[77:60]; // @[EmbeddedTLB.scala 218:70]
  wire [15:0] hitMeta_asid = _T_198[93:78]; // @[EmbeddedTLB.scala 218:70]
  wire [31:0] hitData_pteaddr = _T_198[31:0]; // @[EmbeddedTLB.scala 219:70]
  wire [19:0] hitData_ppn = _T_198[51:32]; // @[EmbeddedTLB.scala 219:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 220:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 220:38]
  reg [2:0] state; // @[EmbeddedTLB.scala 250:22]
  wire  _T_244 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 229:62]
  wire  _T_249 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 229:110]
  wire  _T_251 = ~io_pf_status_sum; // @[EmbeddedTLB.scala 229:137]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u & ~
    io_pf_status_sum); // @[EmbeddedTLB.scala 229:87]
  wire  hitLoad = hitCheck & (hitFlag_r | io_pf_status_mxr & hitFlag_x); // @[EmbeddedTLB.scala 231:26]
  wire  _T_262 = ~io_in_bits_cmd[0] & ~io_in_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_264 = ~hitLoad & _T_262 & hit; // @[EmbeddedTLB.scala 244:40]
  wire  _T_265 = ~ISAMO; // @[EmbeddedTLB.scala 244:50]
  wire  _T_316 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 258:49]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 258:49]
  wire [7:0] _T_307 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,
    memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 295:44]
  reg [1:0] level; // @[EmbeddedTLB.scala 251:22]
  wire  _T_319 = level == 2'h3; // @[EmbeddedTLB.scala 300:58]
  wire  _T_320 = level == 2'h2; // @[EmbeddedTLB.scala 300:73]
  wire  _T_333 = _T_262 & _T_265; // @[EmbeddedTLB.scala 305:38]
  wire  _GEN_19 = ~_T_307[0] | ~_T_307[1] & _T_307[2] ? _T_262 & _T_265 : ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12 301:60 305:22]
  wire  _T_374 = _T_307[0] & ~(_T_244 & ~_T_307[4]) & ~(_T_249 & _T_307[4] & _T_251); // @[EmbeddedTLB.scala 317:87]
  wire  _T_378 = _T_374 & (_T_307[1] | io_pf_status_mxr & _T_307[3]); // @[EmbeddedTLB.scala 319:36]
  wire  _T_379 = _T_374 & _T_307[2]; // @[EmbeddedTLB.scala 320:37]
  wire  _GEN_23 = ~_T_378 & _T_262 | ~_T_379 & io_in_bits_cmd[0] ? _T_333 : ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12 333:80 335:22]
  wire  _GEN_29 = level != 2'h0 ? _GEN_23 : ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12 316:36]
  wire  _GEN_35 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_29; // @[EmbeddedTLB.scala 300:82]
  wire  _GEN_54 = _T_316 ? _GEN_35 : ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12 296:33]
  wire  _GEN_78 = 3'h2 == state ? _GEN_54 : ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12 272:18]
  wire  _GEN_91 = 3'h1 == state ? ~hitLoad & _T_262 & hit & ~ISAMO : _GEN_78; // @[EmbeddedTLB.scala 244:12 272:18]
  wire  loadPF = 3'h0 == state ? ~hitLoad & _T_262 & hit & ~ISAMO : _GEN_91; // @[EmbeddedTLB.scala 244:12 272:18]
  wire  hitStore = hitCheck & hitFlag_w; // @[EmbeddedTLB.scala 232:27]
  wire  _T_335 = io_in_bits_cmd[0] | ISAMO; // @[EmbeddedTLB.scala 306:40]
  wire  _GEN_20 = ~_T_307[0] | ~_T_307[1] & _T_307[2] ? io_in_bits_cmd[0] | ISAMO : ~hitStore & io_in_bits_cmd[0] & hit
     | _T_264 & ISAMO; // @[EmbeddedTLB.scala 245:13 301:60 306:23]
  wire  _GEN_24 = ~_T_378 & _T_262 | ~_T_379 & io_in_bits_cmd[0] ? _T_335 : ~hitStore & io_in_bits_cmd[0] & hit | _T_264
     & ISAMO; // @[EmbeddedTLB.scala 245:13 333:80 336:23]
  wire  _GEN_30 = level != 2'h0 ? _GEN_24 : ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO; // @[EmbeddedTLB.scala 245:13 316:36]
  wire  _GEN_36 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : _GEN_30; // @[EmbeddedTLB.scala 300:82]
  wire  _GEN_55 = _T_316 ? _GEN_36 : ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO; // @[EmbeddedTLB.scala 245:13 296:33]
  wire  _GEN_79 = 3'h2 == state ? _GEN_55 : ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO; // @[EmbeddedTLB.scala 245:13 272:18]
  wire  _GEN_92 = 3'h1 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO : _GEN_79; // @[EmbeddedTLB.scala 245:13 272:18]
  wire  storePF = 3'h0 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO : _GEN_92; // @[EmbeddedTLB.scala 245:13 272:18]
  wire  _T_237 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 136:23]
  wire  hitWB = hit & (~hitFlag_a | ~hitFlag_d & io_in_bits_cmd[0]) & ~(loadPF | storePF | _T_237); // @[EmbeddedTLB.scala 224:81]
  wire [7:0] _T_241 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[Cat.scala 30:58]
  wire [7:0] _T_242 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 225:79]
  wire [7:0] hitRefillFlag = _T_241 | _T_242; // @[EmbeddedTLB.scala 225:69]
  wire [39:0] _T_243 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 30:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  reg  REG_1; // @[EmbeddedTLB.scala 239:26]
  reg  REG_2; // @[EmbeddedTLB.scala 240:27]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 253:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 255:26]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 258:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 259:18]
  wire  _T_292 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_292 | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  wire [31:0] _T_303 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 30:58]
  wire  _T_305 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [8:0] _T_359 = _T_319 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 314:50]
  wire [31:0] _T_361 = {memRdata_ppn,_T_359,3'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_18 = ~_T_307[0] | ~_T_307[1] & _T_307[2] ? 3'h5 : 3'h1; // @[EmbeddedTLB.scala 301:60 302:73 313:19]
  wire [31:0] _GEN_21 = ~_T_307[0] | ~_T_307[1] & _T_307[2] ? raddr : _T_361; // @[EmbeddedTLB.scala 259:18 301:60 314:19]
  wire  _T_384 = ~_T_307[6] | ~_T_307[7] & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 321:72]
  wire [63:0] _T_386 = {56'h0,io_in_bits_cmd[0],7'h40}; // @[Cat.scala 30:58]
  wire [7:0] _T_389 = {_T_307[7],_T_307[6],_T_307[5],_T_307[4],_T_307[3],_T_307[2],_T_307[1],_T_307[0]}; // @[EmbeddedTLB.scala 323:79]
  wire [7:0] _T_390 = _T_241 | _T_389; // @[EmbeddedTLB.scala 323:68]
  wire [63:0] _T_391 = io_mem_resp_bits_rdata | _T_386; // @[EmbeddedTLB.scala 324:50]
  wire [2:0] _T_412 = _T_384 ? 3'h3 : 3'h4; // @[EmbeddedTLB.scala 338:27]
  wire [2:0] _GEN_22 = ~_T_378 & _T_262 | ~_T_379 & io_in_bits_cmd[0] ? 3'h5 : _T_412; // @[EmbeddedTLB.scala 333:80 334:21 338:21]
  wire  _GEN_25 = ~_T_378 & _T_262 | ~_T_379 & io_in_bits_cmd[0] ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 333:80 339:30]
  wire [17:0] _T_415 = _T_320 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 342:59]
  wire [17:0] _T_416 = _T_319 ? 18'h0 : _T_415; // @[EmbeddedTLB.scala 342:26]
  wire [7:0] _GEN_26 = level != 2'h0 ? _T_390 : 8'h0; // @[EmbeddedTLB.scala 316:36 323:26]
  wire [63:0] _GEN_27 = level != 2'h0 ? _T_391 : memRespStore; // @[EmbeddedTLB.scala 316:36 324:24 253:25]
  wire [2:0] _GEN_28 = level != 2'h0 ? _GEN_22 : state; // @[EmbeddedTLB.scala 250:22 316:36]
  wire  _GEN_31 = level != 2'h0 & _GEN_25; // @[EmbeddedTLB.scala 316:36]
  wire [17:0] _GEN_32 = level != 2'h0 ? _T_416 : 18'h3ffff; // @[EmbeddedTLB.scala 316:36 342:20]
  wire [17:0] _GEN_41 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_32; // @[EmbeddedTLB.scala 300:82]
  wire [17:0] _GEN_60 = _T_316 ? _GEN_41 : 18'h3ffff; // @[EmbeddedTLB.scala 296:33]
  wire [17:0] _GEN_84 = 3'h2 == state ? _GEN_60 : 18'h3ffff; // @[EmbeddedTLB.scala 272:18]
  wire [17:0] _GEN_97 = 3'h1 == state ? 18'h3ffff : _GEN_84; // @[EmbeddedTLB.scala 272:18]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_97; // @[EmbeddedTLB.scala 272:18]
  wire [17:0] _GEN_33 = level != 2'h0 ? missMask : missMaskStore; // @[EmbeddedTLB.scala 316:36 343:25 255:26]
  wire [2:0] _GEN_34 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_18 : _GEN_28; // @[EmbeddedTLB.scala 300:82]
  wire [31:0] _GEN_37 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_21 : raddr; // @[EmbeddedTLB.scala 259:18 300:82]
  wire [7:0] _GEN_38 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_26; // @[EmbeddedTLB.scala 300:82]
  wire [63:0] _GEN_39 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_27; // @[EmbeddedTLB.scala 253:25 300:82]
  wire  _GEN_40 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_31; // @[EmbeddedTLB.scala 300:82]
  wire [17:0] _GEN_42 = ~(_T_307[1] | _T_307[3]) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_33; // @[EmbeddedTLB.scala 255:26 300:82]
  wire [1:0] _T_418 = level - 2'h1; // @[EmbeddedTLB.scala 345:24]
  wire [2:0] _GEN_52 = _T_316 ? _GEN_34 : state; // @[EmbeddedTLB.scala 250:22 296:33]
  wire [7:0] _GEN_57 = _T_316 ? _GEN_38 : 8'h0; // @[EmbeddedTLB.scala 296:33]
  wire  _GEN_59 = _T_316 & _GEN_40; // @[EmbeddedTLB.scala 296:33]
  wire [1:0] _GEN_62 = _T_316 ? _T_418 : level; // @[EmbeddedTLB.scala 296:33 345:15 251:22]
  wire [2:0] _GEN_63 = _T_305 ? 3'h4 : state; // @[EmbeddedTLB.scala 250:22 353:{38,46}]
  wire [2:0] _GEN_65 = _GEN_2 ? 3'h0 : state; // @[EmbeddedTLB.scala 356:73 357:13 250:22]
  wire  _GEN_67 = _GEN_2 ? 1'h0 : _GEN_2; // @[EmbeddedTLB.scala 356:73 359:22]
  wire [2:0] _GEN_68 = 3'h5 == state ? 3'h0 : state; // @[EmbeddedTLB.scala 272:18 363:13 250:22]
  wire [2:0] _GEN_69 = 3'h4 == state ? _GEN_65 : _GEN_68; // @[EmbeddedTLB.scala 272:18]
  wire  _GEN_71 = 3'h4 == state ? _GEN_67 : _GEN_2; // @[EmbeddedTLB.scala 272:18]
  wire [2:0] _GEN_72 = 3'h3 == state ? _GEN_63 : _GEN_69; // @[EmbeddedTLB.scala 272:18]
  wire  _GEN_75 = 3'h3 == state ? _GEN_2 : _GEN_71; // @[EmbeddedTLB.scala 272:18]
  wire  _GEN_96 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_59; // @[EmbeddedTLB.scala 272:18]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_96; // @[EmbeddedTLB.scala 272:18]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 368:23]
  wire  _T_436 = state == 3'h0; // @[EmbeddedTLB.scala 374:82]
  reg  REG_7; // @[EmbeddedTLB.scala 374:33]
  reg [3:0] REG_8; // @[EmbeddedTLB.scala 375:21]
  reg [3:0] REG_9; // @[EmbeddedTLB.scala 375:60]
  reg [26:0] REG_10; // @[EmbeddedTLB.scala 375:84]
  reg [15:0] REG_11; // @[EmbeddedTLB.scala 376:19]
  reg [17:0] REG_12; // @[EmbeddedTLB.scala 376:72]
  reg [7:0] REG_13; // @[EmbeddedTLB.scala 377:19]
  reg [19:0] REG_14; // @[EmbeddedTLB.scala 377:77]
  reg [31:0] REG_15; // @[EmbeddedTLB.scala 378:22]
  wire [59:0] lo_6 = {REG_13,REG_14,REG_15}; // @[Cat.scala 30:58]
  wire [60:0] hi_13 = {REG_10,REG_11,REG_12}; // @[Cat.scala 30:58]
  wire [31:0] _T_452 = {hitData_ppn,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_454 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_455 = _T_452 & _T_454; // @[BitUtils.scala 32:13]
  wire [31:0] _T_456 = ~_T_454; // @[BitUtils.scala 32:38]
  wire [31:0] _T_457 = io_in_bits_addr[31:0] & _T_456; // @[BitUtils.scala 32:36]
  wire [31:0] _T_458 = _T_455 | _T_457; // @[BitUtils.scala 32:25]
  wire [31:0] _T_471 = {memRespStore[29:10],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_473 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_474 = _T_471 & _T_473; // @[BitUtils.scala 32:13]
  wire [31:0] _T_475 = ~_T_473; // @[BitUtils.scala 32:38]
  wire [31:0] _T_476 = io_in_bits_addr[31:0] & _T_475; // @[BitUtils.scala 32:36]
  wire [31:0] _T_477 = _T_474 | _T_476; // @[BitUtils.scala 32:25]
  wire  _T_479 = ~hitWB; // @[EmbeddedTLB.scala 383:45]
  wire  _T_486 = hit & ~hitWB ? ~(_T_237 | loadPF | storePF) : state == 3'h4; // @[EmbeddedTLB.scala 383:37]
  assign io_in_ready = io_out_ready & _T_436 & ~miss & _T_479 & io_mdReady & (~_T_237 & ~loadPF & ~storePF); // @[EmbeddedTLB.scala 385:86]
  assign io_out_valid = io_in_valid & _T_486; // @[EmbeddedTLB.scala 383:31]
  assign io_out_bits_addr = hit ? _T_458 : _T_477; // @[EmbeddedTLB.scala 382:26]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 381:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 381:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 381:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 381:15]
  assign io_mdWrite_wen = REG_7; // @[TLB.scala 214:14]
  assign io_mdWrite_windex = REG_8; // @[TLB.scala 215:17]
  assign io_mdWrite_waymask = REG_9; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {hi_13,lo_6}; // @[Cat.scala 30:58]
  assign io_mem_req_valid = state == 3'h1 | cmd; // @[EmbeddedTLB.scala 370:48]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 369:35]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[EmbeddedTLB.scala 369:138]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 371:21]
  assign io_pf_loadPF = REG_1; // @[EmbeddedTLB.scala 239:16]
  assign io_pf_storePF = REG_2; // @[EmbeddedTLB.scala 240:17]
  assign io_pf_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 204:11]
  assign io_isFinish = _T_292 | _T_237; // @[EmbeddedTLB.scala 388:32]
  always @(posedge clock) begin
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_185;
    end
    if (reset) begin // @[EmbeddedTLB.scala 250:22]
      state <= 3'h0; // @[EmbeddedTLB.scala 250:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (hitWB) begin // @[EmbeddedTLB.scala 274:32]
        state <= 3'h3; // @[EmbeddedTLB.scala 275:15]
      end else if (miss) begin // @[EmbeddedTLB.scala 278:37]
        state <= 3'h1; // @[EmbeddedTLB.scala 279:15]
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (_T_305) begin // @[EmbeddedTLB.scala 291:38]
        state <= 3'h2; // @[EmbeddedTLB.scala 291:46]
      end
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      state <= _GEN_52;
    end else begin
      state <= _GEN_72;
    end
    if (reset) begin // @[EmbeddedTLB.scala 251:22]
      level <= 2'h3; // @[EmbeddedTLB.scala 251:22]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (!(hitWB)) begin // @[EmbeddedTLB.scala 274:32]
        if (miss) begin // @[EmbeddedTLB.scala 278:37]
          level <= 2'h3; // @[EmbeddedTLB.scala 281:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
        level <= _GEN_62;
      end
    end
    if (hitWB) begin // @[Reg.scala 16:19]
      hitWBStore <= _T_243; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 239:26]
      REG_1 <= 1'h0; // @[EmbeddedTLB.scala 239:26]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_1 <= ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12]
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_1 <= ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12]
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_1 <= _GEN_54;
    end else begin
      REG_1 <= ~hitLoad & _T_262 & hit & ~ISAMO; // @[EmbeddedTLB.scala 244:12]
    end
    if (reset) begin // @[EmbeddedTLB.scala 240:27]
      REG_2 <= 1'h0; // @[EmbeddedTLB.scala 240:27]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_2 <= ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO; // @[EmbeddedTLB.scala 245:13]
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_2 <= ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO; // @[EmbeddedTLB.scala 245:13]
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_2 <= _GEN_55;
    end else begin
      REG_2 <= ~hitStore & io_in_bits_cmd[0] & hit | _T_264 & ISAMO; // @[EmbeddedTLB.scala 245:13]
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
          if (_T_316) begin // @[EmbeddedTLB.scala 296:33]
            memRespStore <= _GEN_39;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
        if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
          if (_T_316) begin // @[EmbeddedTLB.scala 296:33]
            missMaskStore <= _GEN_42;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (!(hitWB)) begin // @[EmbeddedTLB.scala 274:32]
        if (miss) begin // @[EmbeddedTLB.scala 278:37]
          raddr <= _T_303; // @[EmbeddedTLB.scala 280:15]
        end
      end
    end else if (!(3'h1 == state)) begin // @[EmbeddedTLB.scala 272:18]
      if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
        if (_T_316) begin // @[EmbeddedTLB.scala 296:33]
          raddr <= _GEN_37;
        end
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      if (hitWB) begin // @[EmbeddedTLB.scala 274:32]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 277:24]
      end else if (miss) begin // @[EmbeddedTLB.scala 278:37]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 283:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_75;
    end
    if (reset) begin // @[EmbeddedTLB.scala 374:33]
      REG_7 <= 1'h0; // @[EmbeddedTLB.scala 374:33]
    end else begin
      REG_7 <= missMetaRefill | hitWB & state == 3'h0; // @[EmbeddedTLB.scala 374:33]
    end
    REG_8 <= io_in_bits_addr[15:12]; // @[TLB.scala 200:19]
    if (hit) begin // @[EmbeddedTLB.scala 212:20]
      REG_9 <= hitVec;
    end else begin
      REG_9 <= victimWaymask;
    end
    REG_10 <= {hi,vpn_vpn0}; // @[EmbeddedTLB.scala 375:89]
    if (hitWB) begin // @[EmbeddedTLB.scala 376:23]
      REG_11 <= hitMeta_asid;
    end else begin
      REG_11 <= satp_asid;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 376:76]
      REG_12 <= hitMeta_mask;
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_12 <= 18'h3ffff;
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_12 <= 18'h3ffff;
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_12 <= _GEN_60;
    end else begin
      REG_12 <= 18'h3ffff;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 377:23]
      REG_13 <= hitRefillFlag;
    end else if (3'h0 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_13 <= 8'h0;
    end else if (3'h1 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_13 <= 8'h0;
    end else if (3'h2 == state) begin // @[EmbeddedTLB.scala 272:18]
      REG_13 <= _GEN_57;
    end else begin
      REG_13 <= 8'h0;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 377:81]
      REG_14 <= hitData_ppn;
    end else begin
      REG_14 <= memRdata_ppn;
    end
    if (hitWB) begin // @[EmbeddedTLB.scala 378:27]
      REG_15 <= hitData_pteaddr;
    end else begin
      REG_15 <= raddr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  hitWBStore = _RAND_3[39:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_2 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  memRespStore = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  missMaskStore = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  raddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  alreadyOutFire = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_8 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  REG_9 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  REG_10 = _RAND_13[26:0];
  _RAND_14 = {1{`RANDOM}};
  REG_11 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  REG_12 = _RAND_15[17:0];
  _RAND_16 = {1{`RANDOM}};
  REG_13 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  REG_14 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  REG_15 = _RAND_18[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBEmpty_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  assign io_in_ready = io_out_ready; // @[EmbeddedTLB.scala 406:10]
  assign io_out_valid = io_in_valid; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 406:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 406:10]
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_windex,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  input  [3:0]   io_rindex,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_0_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_0_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_0_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_1 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_1_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_1_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_1_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_2 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_2_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_2_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_2_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg [120:0] tlbmd_3 [0:15]; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_en; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_3_MPORT_addr; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 51:18]
  wire [120:0] tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
  wire [3:0] tlbmd_3_MPORT_1_addr; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_mask; // @[EmbeddedTLB.scala 51:18]
  wire  tlbmd_3_MPORT_1_en; // @[EmbeddedTLB.scala 51:18]
  reg  resetState; // @[EmbeddedTLB.scala 55:27]
  reg [3:0] resetSet; // @[Counter.scala 60:40]
  wire  wrap_wrap = resetSet == 4'hf; // @[Counter.scala 72:24]
  wire [3:0] _wrap_value_T_1 = resetSet + 4'h1; // @[Counter.scala 76:24]
  wire  resetFinish = resetState & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[EmbeddedTLB.scala 57:22 55:27 57:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 66:20]
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = io_rindex;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = io_rindex;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = io_rindex;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = io_rindex;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[EmbeddedTLB.scala 51:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 52:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 72:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 51:18]
    end
    resetState <= reset | _GEN_2; // @[EmbeddedTLB.scala 55:{27,27}]
    if (reset) begin // @[Counter.scala 60:40]
      resetSet <= 4'h0; // @[Counter.scala 60:40]
    end else if (resetState) begin // @[Counter.scala 118:17]
      resetSet <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_csrMMU_status_sum,
  input         io_csrMMU_status_mxr,
  output        io_csrMMU_loadPF,
  output        io_csrMMU_storePF,
  output [38:0] io_csrMMU_addr,
  output        _T_28_0,
  input  [63:0] CSRSATP,
  input         amoReq,
  output        vmEnable_0,
  output        _T_27_0,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 83:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 83:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[EmbeddedTLB.scala 83:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[EmbeddedTLB.scala 83:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 83:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 83:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 83:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[EmbeddedTLB.scala 83:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 83:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 83:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 83:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 83:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 83:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 83:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 83:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_pf_status_sum; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_pf_status_mxr; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 83:23]
  wire [38:0] tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 83:23]
  wire  tlbExec_ISAMO; // @[EmbeddedTLB.scala 83:23]
  wire  tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 84:24]
  wire  tlbEmpty_io_in_valid; // @[EmbeddedTLB.scala 84:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[EmbeddedTLB.scala 84:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[EmbeddedTLB.scala 84:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[EmbeddedTLB.scala 84:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[EmbeddedTLB.scala 84:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[EmbeddedTLB.scala 84:24]
  wire  tlbEmpty_io_out_ready; // @[EmbeddedTLB.scala 84:24]
  wire  tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 84:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 84:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 84:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 84:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 84:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 84:24]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 85:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 85:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 85:21]
  wire [3:0] mdTLB_io_write_windex; // @[EmbeddedTLB.scala 85:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 85:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 85:21]
  wire [3:0] mdTLB_io_rindex; // @[EmbeddedTLB.scala 85:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 85:21]
  reg [120:0] r__0; // @[Reg.scala 15:16]
  reg [120:0] r__1; // @[Reg.scala 15:16]
  reg [120:0] r__2; // @[Reg.scala 15:16]
  reg [120:0] r__3; // @[Reg.scala 15:16]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 117:26]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 105:57]
  reg  REG; // @[EmbeddedTLB.scala 108:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : REG; // @[EmbeddedTLB.scala 108:24 109:{25,33}]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[EmbeddedTLB.scala 110:{50,58}]
  reg [38:0] r_1_addr; // @[Reg.scala 15:16]
  reg [2:0] r_1_size; // @[Reg.scala 15:16]
  reg [3:0] r_1_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_1_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_1_wdata; // @[Reg.scala 15:16]
  wire  _T_15 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_12 = _T_15 ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_16 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_13 = tlbExec_io_out_valid & tlbEmpty_io_in_ready | _GEN_12; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_2_addr; // @[Reg.scala 15:16]
  reg [2:0] r_2_size; // @[Reg.scala 15:16]
  reg [3:0] r_2_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_2_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_2_wdata; // @[Reg.scala 15:16]
  wire  _T_21 = tlbExec_io_out_valid & ~tlbExec_io_out_ready; // @[EmbeddedTLB.scala 145:81]
  reg  r_3; // @[Reg.scala 27:20]
  wire  _GEN_29 = _T_21 | r_3; // @[Reg.scala 28:19 27:20 28:23]
  wire  _T_22 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_26 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[Bundle.scala 136:23]
  wire  _T_27 = tlbExec_io_out_valid & ~r_3 | _T_26; // @[EmbeddedTLB.scala 147:65]
  wire  _T_28 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[Bundle.scala 136:23]
  EmbeddedTLBExec_1 tlbExec ( // @[EmbeddedTLB.scala 83:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_addr(tlbExec_io_pf_addr),
    .io_isFinish(tlbExec_io_isFinish),
    .ISAMO(tlbExec_ISAMO)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[EmbeddedTLB.scala 84:24]
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[EmbeddedTLB.scala 85:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 113:16 126:19 130:21]
  assign io_in_resp_valid = io_out_resp_valid; // @[EmbeddedTLB.scala 141:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 141:15]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 126:19 129:22 138:41]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 126:19 131:26 138:41]
  assign io_out_req_bits_size = ~vmEnable ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 126:19 132:26 138:41]
  assign io_out_req_bits_cmd = ~vmEnable ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 126:19 133:25 138:41]
  assign io_out_req_bits_wmask = ~vmEnable ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 126:19 134:27 138:41]
  assign io_out_req_bits_wdata = ~vmEnable ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 126:19 135:27 138:41]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 90:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 90:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 90:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 90:18]
  assign io_csrMMU_loadPF = tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 91:17]
  assign io_csrMMU_storePF = tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 91:17]
  assign io_csrMMU_addr = tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 91:17]
  assign _T_28_0 = _T_28;
  assign vmEnable_0 = vmEnable;
  assign _T_27_0 = _T_27;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = REG; // @[EmbeddedTLB.scala 115:17]
  assign tlbExec_io_in_bits_addr = r_1_addr; // @[EmbeddedTLB.scala 114:16]
  assign tlbExec_io_in_bits_size = r_1_size; // @[EmbeddedTLB.scala 114:16]
  assign tlbExec_io_in_bits_cmd = r_1_cmd; // @[EmbeddedTLB.scala 114:16]
  assign tlbExec_io_in_bits_wmask = r_1_wmask; // @[EmbeddedTLB.scala 114:16]
  assign tlbExec_io_in_bits_wdata = r_1_wdata; // @[EmbeddedTLB.scala 114:16]
  assign tlbExec_io_out_ready = ~vmEnable | tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 126:19 127:26 Pipeline.scala 29:16]
  assign tlbExec_io_md_0 = r__0; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_md_1 = r__1; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_md_2 = r__2; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_md_3 = r__3; // @[EmbeddedTLB.scala 92:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 93:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 90:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 90:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 90:18]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 89:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 91:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[EmbeddedTLB.scala 91:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 91:17]
  assign tlbExec_ISAMO = amoReq;
  assign tlbEmpty_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = r_2_addr; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = r_2_size; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = r_2_cmd; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = r_2_wmask; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = r_2_wdata; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = ~vmEnable | io_out_req_ready; // @[EmbeddedTLB.scala 126:19 128:52 138:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 102:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 95:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 95:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 95:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 95:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[TLB.scala 200:19]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__0 <= mdTLB_io_tlbmd_0; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__1 <= mdTLB_io_tlbmd_1; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__2 <= mdTLB_io_tlbmd_2; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r__3 <= mdTLB_io_tlbmd_3; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 108:24]
      REG <= 1'h0; // @[EmbeddedTLB.scala 108:24]
    end else begin
      REG <= _GEN_5;
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r_1_addr <= io_in_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r_1_size <= io_in_req_bits_size; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r_1_cmd <= io_in_req_bits_cmd; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r_1_wmask <= io_in_req_bits_wmask; // @[Reg.scala 16:23]
    end
    if (mdUpdate) begin // @[Reg.scala 16:19]
      r_1_wdata <= io_in_req_bits_wdata; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG_1 <= _GEN_13;
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      r_2_addr <= tlbExec_io_out_bits_addr; // @[Reg.scala 16:23]
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      r_2_size <= tlbExec_io_out_bits_size; // @[Reg.scala 16:23]
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      r_2_cmd <= tlbExec_io_out_bits_cmd; // @[Reg.scala 16:23]
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      r_2_wmask <= tlbExec_io_out_bits_wmask; // @[Reg.scala 16:23]
    end
    if (_T_16) begin // @[Reg.scala 16:19]
      r_2_wdata <= tlbExec_io_out_bits_wdata; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3 <= 1'h0; // @[Reg.scala 27:20]
    end else if (r_3 & _T_22) begin // @[EmbeddedTLB.scala 146:53]
      r_3 <= 1'h0; // @[EmbeddedTLB.scala 146:72]
    end else begin
      r_3 <= _GEN_29;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  r__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  r__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  r__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  r__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  r_1_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_size = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  r_1_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  r_1_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  REG_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_2_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  r_2_size = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  r_2_cmd = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  r_2_wmask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  r_2_wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  r_3 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_16 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_16) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 147:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 146:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 145:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 145:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 145:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 145:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 145:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module CacheStage2_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [18:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_dirty,
  output [18:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_dirty,
  output [18:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_dirty,
  output [18:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 176:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 176:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 176:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 178:64]
  reg  isForwardMetaReg; // @[Cache.scala 179:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 180:24 179:33 180:43]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 181:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 181:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 15:16 16:{19,23}]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 15:16 16:{19,23}]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 15:16 16:{19,23}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 185:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 187:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 187:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 187:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 187:61]
  wire [18:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[Cache.scala 189:22]
  wire [18:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[Cache.scala 189:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 192:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_39 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_42 = {_T_39,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 193:42]
  wire  _T_45 = ~metaWay_0_valid; // @[Cache.scala 195:45]
  wire  _T_46 = ~metaWay_1_valid; // @[Cache.scala 195:45]
  wire  _T_47 = ~metaWay_2_valid; // @[Cache.scala 195:45]
  wire  _T_48 = ~metaWay_3_valid; // @[Cache.scala 195:45]
  wire [3:0] invalidVec = {_T_48,_T_47,_T_46,_T_45}; // @[Cache.scala 195:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 196:34]
  wire [1:0] _T_52 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 199:8]
  wire [2:0] _T_53 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_52}; // @[Cache.scala 198:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_53}; // @[Cache.scala 197:33]
  wire [3:0] _T_54 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 202:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  wire [1:0] _T_59 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_61 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_63 = _T_59 + _T_61; // @[Bitwise.scala 47:55]
  wire  _T_65 = _T_63 > 3'h1; // @[Cache.scala 203:26]
  wire [31:0] _T_172 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 87:11]
  wire  _T_174 = _T_172[31:28] == 4'h0; // @[NutCore.scala 87:44]
  wire [31:0] _T_175 = io_in_bits_req_addr ^ 32'h40600000; // @[NutCore.scala 87:11]
  wire  _T_177 = _T_175[31:24] == 8'h0; // @[NutCore.scala 87:44]
  wire [9:0] _T_187 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_189 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_187; // @[Cache.scala 219:13]
  wire  isForwardData = io_in_valid & _T_189; // @[Cache.scala 218:35]
  reg  isForwardDataReg; // @[Cache.scala 221:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 222:24 221:33 222:43]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_196 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_196; // @[Cache.scala 230:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 229:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 228:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 228:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 228:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 228:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 228:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 215:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 213:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  assign io_out_bits_mmio = _T_174 | _T_177; // @[NutCore.scala 88:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 225:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 226:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 226:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 179:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 179:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 181:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 181:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_42;
    end
    if (reset) begin // @[Cache.scala 221:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 221:33]
    end else if (_T_12) begin // @[Cache.scala 223:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 223:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 16:23]
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:210 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 210:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fatal; // @[Cache.scala 210:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  REG = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage3_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [18:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_dirty,
  input  [18:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_dirty,
  input  [18:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_dirty,
  input  [18:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid,
  output [3:0]  io_cohResp_bits_cmd,
  output [63:0] io_cohResp_bits_rdata,
  output        io_dataReadRespToL1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 256:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 256:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 256:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 256:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 256:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 256:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 256:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 257:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 257:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 257:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 257:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 260:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 260:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 261:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 262:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 263:26]
  wire  _T_6 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_6; // @[Cache.scala 264:39]
  wire  _T_7 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_7; // @[Cache.scala 265:26]
  wire  meta_dirty = io_in_bits_waymask[0] & io_in_bits_metas_0_dirty | io_in_bits_waymask[1] & io_in_bits_metas_1_dirty
     | io_in_bits_waymask[2] & io_in_bits_metas_2_dirty | io_in_bits_waymask[3] & io_in_bits_metas_3_dirty; // @[Mux.scala 27:72]
  wire [18:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [18:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 275:49]
  wire [63:0] _T_43 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_43 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_48 | _T_46; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_49; // @[Cache.scala 277:21]
  wire [7:0] _T_62 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_64 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_66 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_77 = {_T_76,_T_74,_T_72,_T_70,_T_68,_T_66,_T_64,_T_62}; // @[Cat.scala 30:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_77 : 64'h0; // @[Cache.scala 278:21]
  reg [2:0] value; // @[Counter.scala 60:40]
  wire  _T_78 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_79 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 281:34]
  wire  _T_80 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_81 = io_in_bits_req_cmd == 4'h3 | _T_80; // @[Cache.scala 281:62]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_0 = _T_78 & (io_in_bits_req_cmd == 4'h3 | _T_80) ? _value_T_1 : value; // @[Cache.scala 281:85 Counter.scala 76:15 60:40]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 285:22]
  wire [63:0] _T_84 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_85 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_86 = dataRead & _T_85; // @[BitUtils.scala 32:36]
  wire [2:0] _T_91 = _T_81 ? value : addr_wordIndex; // @[Cache.scala 288:51]
  wire  metaHitWriteBus_req_valid = hitWrite & ~meta_dirty; // @[Cache.scala 291:22]
  reg [3:0] state; // @[Cache.scala 296:22]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 306:23]
  wire  _T_103 = state == 4'h3; // @[Cache.scala 308:39]
  wire  _T_104 = state == 4'h8; // @[Cache.scala 308:66]
  wire [2:0] _T_109 = _T_104 ? value_1 : value_2; // @[Cache.scala 309:33]
  wire  _T_111 = state2 == 2'h1; // @[Cache.scala 310:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_116 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_117 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_118 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_119 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_120 = _T_116 | _T_117; // @[Mux.scala 27:72]
  wire [63:0] _T_121 = _T_120 | _T_118; // @[Mux.scala 27:72]
  wire  _T_124 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_127 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_130 = hitReadBurst & io_out_ready; // @[Cache.scala 316:83]
  wire [1:0] _GEN_8 = _T_127 | io_cohResp_valid | hitReadBurst & io_out_ready ? 2'h0 : state2; // @[Cache.scala 316:{100,109} 306:23]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_133 = state == 4'h1; // @[Cache.scala 324:23]
  wire [2:0] _T_135 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 325:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_135; // @[Cache.scala 324:16]
  wire  _T_141 = state2 == 2'h2; // @[Cache.scala 331:89]
  reg  afterFirstRead; // @[Cache.scala 338:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_78 | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  wire  _T_147 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_149 = state == 4'h2; // @[Cache.scala 340:70]
  wire  readingFirst = ~afterFirstRead & _T_147 & state == 4'h2; // @[Cache.scala 340:60]
  wire  _T_152 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 342:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_153 = state == 4'h0; // @[Cache.scala 345:31]
  wire  _T_157 = _T_104 & _T_141; // @[Cache.scala 346:46]
  wire  _T_161 = _T_104 & io_cohResp_valid; // @[Cache.scala 348:49]
  reg [2:0] value_3; // @[Counter.scala 60:40]
  wire  wrap_wrap = value_3 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_1 = value_3 + 3'h1; // @[Counter.scala 76:24]
  wire  releaseLast = _T_161 & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire [2:0] _T_163 = releaseLast ? 3'h6 : 3'h0; // @[Cache.scala 349:54]
  wire [3:0] _T_164 = hit ? 4'hc : 4'h8; // @[Cache.scala 350:8]
  wire  respToL1Fire = _T_130 & _T_141; // @[Cache.scala 352:51]
  wire  _T_174 = (_T_153 | _T_157) & hitReadBurst & io_out_ready; // @[Cache.scala 353:112]
  reg [2:0] value_4; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = value_4 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_3 = value_4 + 3'h1; // @[Counter.scala 76:24]
  wire  respToL1Last = _T_174 & wrap_wrap_1; // @[Counter.scala 118:{17,24}]
  wire [3:0] _T_177 = hit ? 4'h8 : 4'h0; // @[Cache.scala 362:23]
  wire [2:0] _value_T_4 = addr_wordIndex + 3'h1; // @[Cache.scala 367:93]
  wire [2:0] _value_T_5 = addr_wordIndex == 3'h7 ? 3'h0 : _value_T_4; // @[Cache.scala 367:33]
  wire [3:0] _T_184 = meta_dirty ? 4'h3 : 4'h1; // @[Cache.scala 369:42]
  wire [3:0] _T_185 = mmio ? 4'h5 : _T_184; // @[Cache.scala 369:21]
  wire [3:0] _GEN_20 = miss | mmio ? _T_185 : state; // @[Cache.scala 368:49 369:15 296:22]
  wire  _T_187 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_189 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = _T_189 ? 4'h7 : state; // @[Cache.scala 296:22 374:{50,58}]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid | respToL1Fire ? _value_T_7 : value_1; // @[Cache.scala 377:48 Counter.scala 76:15 60:40]
  wire [3:0] _GEN_28 = probe & io_cohResp_valid & releaseLast | respToL1Fire & respToL1Last ? 4'h0 : state; // @[Cache.scala 296:22 378:{88,96}]
  wire [3:0] _GEN_29 = _T_127 ? 4'h2 : state; // @[Cache.scala 381:50 382:13 296:22]
  wire [2:0] _GEN_30 = _T_127 ? addr_wordIndex : value_1; // @[Cache.scala 381:50 383:25 Counter.scala 60:40]
  wire [2:0] _GEN_31 = _T_79 ? 3'h0 : _GEN_0; // @[Cache.scala 390:{52,75}]
  wire  _T_203 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_203 ? 4'h7 : state; // @[Cache.scala 296:22 391:{46,54}]
  wire  _GEN_33 = _T_147 | afterFirstRead; // @[Cache.scala 387:33 388:24 338:31]
  wire [2:0] _GEN_34 = _T_147 ? _value_T_7 : value_1; // @[Cache.scala 387:33 Counter.scala 76:15 60:40]
  wire [2:0] _GEN_35 = _T_147 ? _GEN_31 : _GEN_0; // @[Cache.scala 387:33]
  wire [3:0] _GEN_36 = _T_147 ? _GEN_32 : state; // @[Cache.scala 296:22 387:33]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_127 ? _value_T_11 : value_2; // @[Cache.scala 396:32 Counter.scala 76:15 60:40]
  wire  _T_206 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_206 & _T_127 ? 4'h4 : state; // @[Cache.scala 296:22 397:{65,73}]
  wire [3:0] _GEN_39 = _T_147 ? 4'h1 : state; // @[Cache.scala 296:22 400:{53,61}]
  wire [3:0] _GEN_40 = _GEN_12 ? 4'h0 : state; // @[Cache.scala 296:22 401:{76,84}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[Cache.scala 355:18 296:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[Cache.scala 355:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : value_2; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[Cache.scala 355:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : value_1; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [2:0] _GEN_47 = 4'h2 == state ? _GEN_35 : _GEN_0; // @[Cache.scala 355:18]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[Cache.scala 355:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? value_2 : _GEN_43; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[Cache.scala 355:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[Cache.scala 355:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_53 = 4'h1 == state ? _GEN_0 : _GEN_47; // @[Cache.scala 355:18]
  wire [2:0] _GEN_54 = 4'h1 == state ? value_2 : _GEN_49; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[Cache.scala 355:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? _GEN_28 : _GEN_50; // @[Cache.scala 355:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_58 = 4'h8 == state ? _GEN_0 : _GEN_53; // @[Cache.scala 355:18]
  wire [2:0] _GEN_59 = 4'h8 == state ? value_2 : _GEN_54; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [63:0] _T_215 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 404:67]
  wire [63:0] _T_216 = io_in_bits_req_wdata & _T_215; // @[BitUtils.scala 32:13]
  wire [63:0] _T_217 = ~_T_215; // @[BitUtils.scala 32:38]
  wire [63:0] _T_218 = io_mem_resp_bits_rdata & _T_217; // @[BitUtils.scala 32:36]
  wire  dataRefillWriteBus_req_valid = _T_149 & _T_147; // @[Cache.scala 406:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_203; // @[Cache.scala 414:61]
  wire  _T_240 = ~io_in_bits_req_cmd[0] & ~io_in_bits_req_cmd[3]; // @[SimpleBus.scala 73:26]
  wire [2:0] _T_242 = io_in_bits_req_cmd[0] ? 3'h5 : 3'h0; // @[Cache.scala 442:79]
  wire [2:0] _T_243 = _T_240 ? 3'h6 : _T_242; // @[Cache.scala 442:27]
  wire  _T_248 = state == 4'h7; // @[Cache.scala 448:48]
  wire  _T_267 = io_in_bits_req_cmd[0] | mmio ? _T_248 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 449:45]
  wire  _T_269 = probe ? 1'h0 : hit | _T_267; // @[Cache.scala 449:8]
  wire  _T_276 = miss ? _T_153 : _T_104 & releaseLast; // @[Cache.scala 456:53]
  wire  _T_285 = hit | io_in_bits_req_cmd[0] ? _T_78 : _T_248 & _GEN_12; // @[Cache.scala 457:8]
  Arbiter metaWriteArb ( // @[Cache.scala 256:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 257:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & (_T_153 & ~hitReadBurst) & ~miss & ~probe; // @[Cache.scala 460:79]
  assign io_out_valid = io_in_valid & _T_269; // @[Cache.scala 447:31]
  assign io_out_bits_cmd = {{1'd0}, _T_243}; // @[Cache.scala 442:21]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 441:29]
  assign io_isFinish = probe ? io_cohResp_valid & _T_276 : _T_285; // @[Cache.scala 456:21]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 308:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_109}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 411:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 421:23]
  assign io_mem_req_valid = _T_133 | _T_103 & state2 == 2'h2; // @[Cache.scala 331:48]
  assign io_mem_req_bits_addr = _T_133 ? raddr : waddr; // @[Cache.scala 326:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_121 | _T_119; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 330:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 336:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 334:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[Cache.scala 334:20]
  assign io_mmio_req_bits_cmd = io_in_bits_req_cmd; // @[Cache.scala 334:20]
  assign io_mmio_req_bits_wmask = io_in_bits_req_wmask; // @[Cache.scala 334:20]
  assign io_mmio_req_bits_wdata = io_in_bits_req_wdata; // @[Cache.scala 334:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 335:22]
  assign io_cohResp_valid = state == 4'h0 & probe | _T_157; // @[Cache.scala 345:53]
  assign io_cohResp_bits_cmd = _T_104 ? {{1'd0}, _T_163} : _T_164; // @[Cache.scala 349:29]
  assign io_cohResp_bits_rdata = _T_121 | _T_119; // @[Mux.scala 27:72]
  assign io_dataReadRespToL1 = hitReadBurst & (_T_153 & io_out_ready | _T_157); // @[Cache.scala 461:39]
  assign metaWriteArb_io_in_0_valid = hitWrite & ~meta_dirty; // @[Cache.scala 291:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h1; // @[Cache.scala 292:16 97:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 290:29 SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_203; // @[Cache.scala 414:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 260:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[SimpleBus.scala 74:22]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 413:32 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 285:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_91}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = _T_84 | _T_86; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 286:29 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _T_149 & _T_147; // @[Cache.scala 406:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = _T_216 | _T_218; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:32 SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      value <= _GEN_0;
    end else if (4'h5 == state) begin // @[Cache.scala 355:18]
      value <= _GEN_0;
    end else if (4'h6 == state) begin // @[Cache.scala 355:18]
      value <= _GEN_0;
    end else begin
      value <= _GEN_58;
    end
    if (reset) begin // @[Cache.scala 296:22]
      state <= 4'h0; // @[Cache.scala 296:22]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      if (probe) begin // @[Cache.scala 360:20]
        if (io_cohResp_valid) begin // @[Cache.scala 361:34]
          state <= _T_177; // @[Cache.scala 362:17]
        end
      end else if (_T_130) begin // @[Cache.scala 365:50]
        state <= 4'h8; // @[Cache.scala 366:15]
      end else begin
        state <= _GEN_20;
      end
    end else if (4'h5 == state) begin // @[Cache.scala 355:18]
      if (_T_187) begin // @[Cache.scala 373:48]
        state <= 4'h6; // @[Cache.scala 373:56]
      end
    end else if (4'h6 == state) begin // @[Cache.scala 355:18]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      if (probe) begin // @[Cache.scala 360:20]
        if (io_cohResp_valid) begin // @[Cache.scala 361:34]
          value_1 <= addr_wordIndex; // @[Cache.scala 363:29]
        end
      end else if (_T_130) begin // @[Cache.scala 365:50]
        value_1 <= _value_T_5; // @[Cache.scala 367:27]
      end
    end else if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
        value_1 <= _GEN_55;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 306:23]
      state2 <= 2'h0; // @[Cache.scala 306:23]
    end else if (2'h0 == state2) begin // @[Cache.scala 313:19]
      if (_T_124) begin // @[Cache.scala 314:53]
        state2 <= 2'h1; // @[Cache.scala 314:62]
      end
    end else if (2'h1 == state2) begin // @[Cache.scala 313:19]
      state2 <= 2'h2; // @[Cache.scala 315:35]
    end else if (2'h2 == state2) begin // @[Cache.scala 313:19]
      state2 <= _GEN_8;
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Cache.scala 338:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 338:31]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      afterFirstRead <= 1'h0; // @[Cache.scala 357:22]
    end else if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      alreadyOutFire <= 1'h0; // @[Cache.scala 358:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_152) begin // @[Reg.scala 16:19]
      if (mmio) begin // @[Cache.scala 341:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_3 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_161) begin // @[Counter.scala 118:17]
      value_3 <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_4 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_174) begin // @[Counter.scala 118:17]
      value_4 <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:267 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 267:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 267:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:463 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 463:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 463:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:464 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 464:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 464:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  value_3 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  value_4 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_9(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_size = io_in_0_valid ? io_in_0_bits_size : io_in_1_bits_size; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_cmd = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_wmask = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : io_in_1_bits_wdata; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module Cache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  output        io_out_coh_req_ready,
  input         io_out_coh_req_valid,
  input  [31:0] io_out_coh_req_bits_addr,
  input  [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_valid,
  output [3:0]  io_out_coh_resp_bits_cmd,
  output [63:0] io_out_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 482:18]
  wire  s1_io_in_valid; // @[Cache.scala 482:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 482:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 482:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 482:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 482:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 482:18]
  wire  s1_io_out_ready; // @[Cache.scala 482:18]
  wire  s1_io_out_valid; // @[Cache.scala 482:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 482:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 482:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 482:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 482:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 482:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 482:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 482:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 482:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 482:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 482:18]
  wire  s2_clock; // @[Cache.scala 483:18]
  wire  s2_reset; // @[Cache.scala 483:18]
  wire  s2_io_in_ready; // @[Cache.scala 483:18]
  wire  s2_io_in_valid; // @[Cache.scala 483:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 483:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 483:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 483:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 483:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 483:18]
  wire  s2_io_out_ready; // @[Cache.scala 483:18]
  wire  s2_io_out_valid; // @[Cache.scala 483:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 483:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 483:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 483:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 483:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 483:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 483:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 483:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 483:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 483:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 483:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 483:18]
  wire  s3_clock; // @[Cache.scala 484:18]
  wire  s3_reset; // @[Cache.scala 484:18]
  wire  s3_io_in_ready; // @[Cache.scala 484:18]
  wire  s3_io_in_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 484:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 484:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 484:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 484:18]
  wire  s3_io_out_ready; // @[Cache.scala 484:18]
  wire  s3_io_out_valid; // @[Cache.scala 484:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_isFinish; // @[Cache.scala 484:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 484:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 484:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 484:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 484:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 484:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 484:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 484:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 484:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 484:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 484:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 484:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 484:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[Cache.scala 484:18]
  wire [3:0] s3_io_mmio_req_bits_cmd; // @[Cache.scala 484:18]
  wire [7:0] s3_io_mmio_req_bits_wmask; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mmio_req_bits_wdata; // @[Cache.scala 484:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 484:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 484:18]
  wire [3:0] s3_io_cohResp_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_cohResp_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 484:18]
  wire  metaArray_clock; // @[Cache.scala 485:25]
  wire  metaArray_reset; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 485:25]
  wire [6:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 485:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 485:25]
  wire [6:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 485:25]
  wire [18:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 485:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 485:25]
  wire  dataArray_clock; // @[Cache.scala 486:25]
  wire  dataArray_reset; // @[Cache.scala 486:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 486:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 486:25]
  wire [9:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 486:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 486:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 486:25]
  wire [9:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 486:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 486:25]
  wire [9:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 486:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 486:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 495:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 495:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 495:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 495:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 495:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 495:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 495:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 495:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 495:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 495:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 495:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 495:19]
  wire  arb_io_out_ready; // @[Cache.scala 495:19]
  wire  arb_io_out_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 495:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 495:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 495:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 495:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 495:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_req_size; // @[Reg.scala 15:16]
  reg [3:0] r_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_req_wdata; // @[Reg.scala 15:16]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_5 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = s2_io_out_valid & s3_io_in_ready | _GEN_8; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [2:0] r_1_req_size; // @[Reg.scala 15:16]
  reg [3:0] r_1_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_1_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_1_req_wdata; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_0_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_0_dirty; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_1_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_1_dirty; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_2_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_2_dirty; // @[Reg.scala 15:16]
  reg [18:0] r_1_metas_3_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_3_data; // @[Reg.scala 15:16]
  reg  r_1_hit; // @[Reg.scala 15:16]
  reg [3:0] r_1_waymask; // @[Reg.scala 15:16]
  reg  r_1_mmio; // @[Reg.scala 15:16]
  reg  r_1_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] r_1_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] r_1_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_11 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  CacheStage1_1 s1 ( // @[Cache.scala 482:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2_1 s2 ( // @[Cache.scala 483:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3_1 s3 ( // @[Cache.scala 484:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(s3_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(s3_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(s3_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_cohResp_bits_cmd(s3_io_cohResp_bits_cmd),
    .io_cohResp_bits_rdata(s3_io_cohResp_bits_rdata),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 485:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 486:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 495:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 496:28]
  assign io_in_resp_valid = s3_io_out_valid & _T_11 ? 1'h0 : s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 512:26]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 506:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 506:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 508:14]
  assign io_out_coh_req_ready = arb_io_in_0_ready; // @[Cache.scala 521:26]
  assign io_out_coh_resp_valid = s3_io_cohResp_valid; // @[Cache.scala 522:21]
  assign io_out_coh_resp_bits_cmd = s3_io_cohResp_bits_cmd; // @[Cache.scala 522:21]
  assign io_out_coh_resp_bits_rdata = s3_io_cohResp_bits_rdata; // @[Cache.scala 522:21]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 509:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 509:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[Cache.scala 509:11]
  assign io_mmio_req_bits_cmd = s3_io_mmio_req_bits_cmd; // @[Cache.scala 509:11]
  assign io_mmio_req_bits_wmask = s3_io_mmio_req_bits_wmask; // @[Cache.scala 509:11]
  assign io_mmio_req_bits_wdata = s3_io_mmio_req_bits_wdata; // @[Cache.scala 509:11]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 498:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 498:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 498:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 498:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 498:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 498:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 530:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 531:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = r_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = r_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = r_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = r_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = r_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 537:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 540:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 539:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = r_1_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = r_1_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = r_1_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = r_1_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = r_1_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = r_1_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = r_1_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = r_1_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = r_1_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = r_1_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = r_1_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = r_1_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = r_1_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = r_1_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = r_1_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = r_1_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = r_1_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = r_1_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = r_1_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = r_1_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = r_1_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = r_1_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = r_1_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 506:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 532:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 508:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 509:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 509:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 509:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 530:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 530:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 534:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 531:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 531:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 532:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 532:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 535:18]
  assign arb_io_in_0_valid = io_out_coh_req_valid; // @[Cache.scala 520:24]
  assign arb_io_in_0_bits_addr = io_out_coh_req_bits_addr; // @[Cache.scala 517:19 SimpleBus.scala 64:15]
  assign arb_io_in_0_bits_size = 3'h3; // @[Cache.scala 517:19 SimpleBus.scala 66:15]
  assign arb_io_in_0_bits_cmd = 4'h8; // @[Cache.scala 517:19 SimpleBus.scala 65:14]
  assign arb_io_in_0_bits_wmask = 8'hff; // @[Cache.scala 517:19 SimpleBus.scala 68:16]
  assign arb_io_in_0_bits_wdata = io_out_coh_req_bits_wdata; // @[Cache.scala 517:19 SimpleBus.scala 67:16]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 496:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 498:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_size <= s1_io_out_bits_req_size; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_cmd <= s1_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wmask <= s1_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wdata <= s1_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG_1 <= _GEN_9;
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_size <= s2_io_out_bits_req_size; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_cmd <= s2_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wmask <= s2_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wdata <= s2_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_hit <= s2_io_out_bits_hit; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  r_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  r_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  r_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_1_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_1_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  r_1_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  r_1_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  r_1_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  r_1_metas_0_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  r_1_metas_0_dirty = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_1_metas_1_tag = _RAND_14[18:0];
  _RAND_15 = {1{`RANDOM}};
  r_1_metas_1_dirty = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_metas_2_tag = _RAND_16[18:0];
  _RAND_17 = {1{`RANDOM}};
  r_1_metas_2_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_1_metas_3_tag = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  r_1_metas_3_dirty = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  r_1_datas_0_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  r_1_datas_1_data = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  r_1_datas_2_data = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  r_1_datas_3_data = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  r_1_hit = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_1_waymask = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  r_1_mmio = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_1_isForwardData = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  r_1_forwardData_data_data = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  r_1_forwardData_waymask = _RAND_29[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready,
  output        io_imem_mem_req_valid,
  output [31:0] io_imem_mem_req_bits_addr,
  output [3:0]  io_imem_mem_req_bits_cmd,
  output [63:0] io_imem_mem_req_bits_wdata,
  input         io_imem_mem_resp_valid,
  input  [3:0]  io_imem_mem_resp_bits_cmd,
  input  [63:0] io_imem_mem_resp_bits_rdata,
  input         io_dmem_mem_req_ready,
  output        io_dmem_mem_req_valid,
  output [31:0] io_dmem_mem_req_bits_addr,
  output [3:0]  io_dmem_mem_req_bits_cmd,
  output [63:0] io_dmem_mem_req_bits_wdata,
  input         io_dmem_mem_resp_valid,
  input  [3:0]  io_dmem_mem_resp_bits_cmd,
  input  [63:0] io_dmem_mem_resp_bits_rdata,
  output        io_dmem_coh_req_ready,
  input         io_dmem_coh_req_valid,
  input  [31:0] io_dmem_coh_req_bits_addr,
  input  [63:0] io_dmem_coh_req_bits_wdata,
  output        io_dmem_coh_resp_valid,
  output [3:0]  io_dmem_coh_resp_bits_cmd,
  output [63:0] io_dmem_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [3:0]  io_mmio_resp_bits_cmd,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_frontend_req_ready,
  input         io_frontend_req_valid,
  input  [31:0] io_frontend_req_bits_addr,
  input  [2:0]  io_frontend_req_bits_size,
  input  [3:0]  io_frontend_req_bits_cmd,
  input  [7:0]  io_frontend_req_bits_wmask,
  input  [63:0] io_frontend_req_bits_wdata,
  input         io_frontend_resp_ready,
  output        io_frontend_resp_valid,
  output [3:0]  io_frontend_resp_bits_cmd,
  output [63:0] io_frontend_resp_bits_rdata,
  output [63:0] perfCnts_2,
  output [38:0] io_in_bits_decode_cf_pc,
  output [4:0]  io_wb_rfDest,
  input         io_extra_mtip,
  input         io_extra_meip_0,
  output        io_wb_rfWen,
  output [63:0] io_wb_rfData,
  input         io_extra_msip,
  output        io_in_valid_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[NutCore.scala 104:34]
  wire  frontend_reset; // @[NutCore.scala 104:34]
  wire  frontend_io_imem_req_ready; // @[NutCore.scala 104:34]
  wire  frontend_io_imem_req_valid; // @[NutCore.scala 104:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[NutCore.scala 104:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[NutCore.scala 104:34]
  wire  frontend_io_imem_resp_ready; // @[NutCore.scala 104:34]
  wire  frontend_io_imem_resp_valid; // @[NutCore.scala 104:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[NutCore.scala 104:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_ready; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_valid; // @[NutCore.scala 104:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[NutCore.scala 104:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[NutCore.scala 104:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_0; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_2; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_4; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_6; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_8; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_10; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[NutCore.scala 104:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 104:34]
  wire [63:0] frontend_io_out_0_bits_cf_runahead_checkpoint_id; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[NutCore.scala 104:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[NutCore.scala 104:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[NutCore.scala 104:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[NutCore.scala 104:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_vtag; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_vec_addr; // @[NutCore.scala 104:34]
  wire [3:0] frontend_io_out_0_bits_ctrl_length_k; // @[NutCore.scala 104:34]
  wire [1:0] frontend_io_out_0_bits_ctrl_algorithm; // @[NutCore.scala 104:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_ready; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_valid; // @[NutCore.scala 104:34]
  wire [63:0] frontend_io_out_1_bits_cf_instr; // @[NutCore.scala 104:34]
  wire [38:0] frontend_io_out_1_bits_cf_pc; // @[NutCore.scala 104:34]
  wire [38:0] frontend_io_out_1_bits_cf_pnpc; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_exceptionVec_1; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_exceptionVec_2; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_exceptionVec_12; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_0; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_1; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_2; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_3; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_4; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_5; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_6; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_7; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_8; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_9; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_10; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_intrVec_11; // @[NutCore.scala 104:34]
  wire [3:0] frontend_io_out_1_bits_cf_brIdx; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_cf_crossPageIPFFix; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_ctrl_src1Type; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_ctrl_src2Type; // @[NutCore.scala 104:34]
  wire [2:0] frontend_io_out_1_bits_ctrl_fuType; // @[NutCore.scala 104:34]
  wire [6:0] frontend_io_out_1_bits_ctrl_fuOpType; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_1_bits_ctrl_rfSrc1; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_1_bits_ctrl_rfSrc2; // @[NutCore.scala 104:34]
  wire  frontend_io_out_1_bits_ctrl_rfWen; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_1_bits_ctrl_rfDest; // @[NutCore.scala 104:34]
  wire [2:0] frontend_io_out_1_bits_ctrl_vtag; // @[NutCore.scala 104:34]
  wire [4:0] frontend_io_out_1_bits_ctrl_vec_addr; // @[NutCore.scala 104:34]
  wire [3:0] frontend_io_out_1_bits_ctrl_length_k; // @[NutCore.scala 104:34]
  wire [1:0] frontend_io_out_1_bits_ctrl_algorithm; // @[NutCore.scala 104:34]
  wire [63:0] frontend_io_out_1_bits_data_imm; // @[NutCore.scala 104:34]
  wire [3:0] frontend_io_flushVec; // @[NutCore.scala 104:34]
  wire [38:0] frontend_io_redirect_target; // @[NutCore.scala 104:34]
  wire  frontend_io_redirect_valid; // @[NutCore.scala 104:34]
  wire  frontend_io_ipf; // @[NutCore.scala 104:34]
  wire  frontend_flushICache; // @[NutCore.scala 104:34]
  wire  frontend_REG_0_valid; // @[NutCore.scala 104:34]
  wire [38:0] frontend_REG_0_pc; // @[NutCore.scala 104:34]
  wire  frontend_REG_0_isMissPredict; // @[NutCore.scala 104:34]
  wire [38:0] frontend_REG_0_actualTarget; // @[NutCore.scala 104:34]
  wire  frontend_REG_0_actualTaken; // @[NutCore.scala 104:34]
  wire [6:0] frontend_REG_0_fuOpType; // @[NutCore.scala 104:34]
  wire [1:0] frontend_REG_0_btbType; // @[NutCore.scala 104:34]
  wire  frontend_REG_0_isRVC; // @[NutCore.scala 104:34]
  wire  frontend_vmEnable; // @[NutCore.scala 104:34]
  wire [11:0] frontend_intrVec; // @[NutCore.scala 104:34]
  wire  frontend_flushTLB; // @[NutCore.scala 104:34]
  wire  Backend_inorder_clock; // @[NutCore.scala 147:25]
  wire  Backend_inorder_reset; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_ready; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_valid; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_io_in_0_bits_cf_instr; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pc; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pnpc; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_1; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_2; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_12; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_0; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_1; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_2; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_3; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_4; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_5; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_6; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_7; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_8; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_9; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_10; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_11; // @[NutCore.scala 147:25]
  wire [3:0] Backend_inorder_io_in_0_bits_cf_brIdx; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_io_in_0_bits_cf_runahead_checkpoint_id; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_src1Type; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_src2Type; // @[NutCore.scala 147:25]
  wire [2:0] Backend_inorder_io_in_0_bits_ctrl_fuType; // @[NutCore.scala 147:25]
  wire [6:0] Backend_inorder_io_in_0_bits_ctrl_fuOpType; // @[NutCore.scala 147:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc1; // @[NutCore.scala 147:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc2; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_rfWen; // @[NutCore.scala 147:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfDest; // @[NutCore.scala 147:25]
  wire [2:0] Backend_inorder_io_in_0_bits_ctrl_vtag; // @[NutCore.scala 147:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_vec_addr; // @[NutCore.scala 147:25]
  wire [3:0] Backend_inorder_io_in_0_bits_ctrl_length_k; // @[NutCore.scala 147:25]
  wire [1:0] Backend_inorder_io_in_0_bits_ctrl_algorithm; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_io_in_0_bits_data_imm; // @[NutCore.scala 147:25]
  wire [1:0] Backend_inorder_io_flush; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_dmem_req_ready; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_dmem_req_valid; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_io_dmem_req_bits_addr; // @[NutCore.scala 147:25]
  wire [2:0] Backend_inorder_io_dmem_req_bits_size; // @[NutCore.scala 147:25]
  wire [3:0] Backend_inorder_io_dmem_req_bits_cmd; // @[NutCore.scala 147:25]
  wire [7:0] Backend_inorder_io_dmem_req_bits_wmask; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_io_dmem_req_bits_wdata; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_dmem_resp_valid; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_io_dmem_resp_bits_rdata; // @[NutCore.scala 147:25]
  wire [1:0] Backend_inorder_io_memMMU_imem_priviledgeMode; // @[NutCore.scala 147:25]
  wire [1:0] Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_memMMU_dmem_status_sum; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_memMMU_dmem_status_mxr; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_memMMU_dmem_loadPF; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_memMMU_dmem_storePF; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_io_memMMU_dmem_addr; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_io_redirect_target; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_redirect_valid; // @[NutCore.scala 147:25]
  wire  Backend_inorder__T_28; // @[NutCore.scala 147:25]
  wire  Backend_inorder_flushICache; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_perfCnts_2; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_io_in_bits_decode_cf_pc; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_satp; // @[NutCore.scala 147:25]
  wire  Backend_inorder_REG_0_valid; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_REG_0_pc; // @[NutCore.scala 147:25]
  wire  Backend_inorder_REG_0_isMissPredict; // @[NutCore.scala 147:25]
  wire [38:0] Backend_inorder_REG_0_actualTarget; // @[NutCore.scala 147:25]
  wire  Backend_inorder_REG_0_actualTaken; // @[NutCore.scala 147:25]
  wire [6:0] Backend_inorder_REG_0_fuOpType; // @[NutCore.scala 147:25]
  wire [1:0] Backend_inorder_REG_0_btbType; // @[NutCore.scala 147:25]
  wire  Backend_inorder_REG_0_isRVC; // @[NutCore.scala 147:25]
  wire [4:0] Backend_inorder_io_wb_rfDest; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_extra_mtip; // @[NutCore.scala 147:25]
  wire  Backend_inorder_amoReq; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_extra_meip_0; // @[NutCore.scala 147:25]
  wire  Backend_inorder_vmEnable; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_wb_rfWen; // @[NutCore.scala 147:25]
  wire [63:0] Backend_inorder_io_wb_rfData; // @[NutCore.scala 147:25]
  wire [11:0] Backend_inorder_intrVec; // @[NutCore.scala 147:25]
  wire  Backend_inorder__T_27; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_extra_msip; // @[NutCore.scala 147:25]
  wire  Backend_inorder_flushTLB; // @[NutCore.scala 147:25]
  wire  Backend_inorder_io_in_valid_0; // @[NutCore.scala 147:25]
  wire  SimpleBusCrossbarNto1_clock; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_reset; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_ready; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_valid; // @[NutCore.scala 151:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_0_req_bits_addr; // @[NutCore.scala 151:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_req_bits_cmd; // @[NutCore.scala 151:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wmask; // @[NutCore.scala 151:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wdata; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[NutCore.scala 151:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd; // @[NutCore.scala 151:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_ready; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_valid; // @[NutCore.scala 151:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_1_req_bits_addr; // @[NutCore.scala 151:26]
  wire [2:0] SimpleBusCrossbarNto1_io_in_1_req_bits_size; // @[NutCore.scala 151:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_req_bits_cmd; // @[NutCore.scala 151:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wmask; // @[NutCore.scala 151:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wdata; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[NutCore.scala 151:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd; // @[NutCore.scala 151:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_out_req_ready; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 151:26]
  wire [31:0] SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 151:26]
  wire [2:0] SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 151:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 151:26]
  wire [7:0] SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 151:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_ready; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_valid; // @[NutCore.scala 151:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_resp_bits_cmd; // @[NutCore.scala 151:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_resp_bits_rdata; // @[NutCore.scala 151:26]
  wire  SimpleBusCrossbarNto1_1_clock; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_reset; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_valid; // @[NutCore.scala 152:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr; // @[NutCore.scala 152:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_size; // @[NutCore.scala 152:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd; // @[NutCore.scala 152:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_valid; // @[NutCore.scala 152:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr; // @[NutCore.scala 152:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_valid; // @[NutCore.scala 152:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr; // @[NutCore.scala 152:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_valid; // @[NutCore.scala 152:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr; // @[NutCore.scala 152:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_size; // @[NutCore.scala 152:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd; // @[NutCore.scala 152:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_ready; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 152:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_ready; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_valid; // @[NutCore.scala 152:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[NutCore.scala 152:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[NutCore.scala 152:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[NutCore.scala 152:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[NutCore.scala 152:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_valid; // @[NutCore.scala 152:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd; // @[NutCore.scala 152:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata; // @[NutCore.scala 152:26]
  wire  EmbeddedTLB_clock; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_reset; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_in_req_valid; // @[EmbeddedTLB.scala 421:23]
  wire [38:0] EmbeddedTLB_io_in_req_bits_addr; // @[EmbeddedTLB.scala 421:23]
  wire [86:0] EmbeddedTLB_io_in_req_bits_user; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_in_resp_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 421:23]
  wire [86:0] EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_out_req_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_out_req_valid; // @[EmbeddedTLB.scala 421:23]
  wire [31:0] EmbeddedTLB_io_out_req_bits_addr; // @[EmbeddedTLB.scala 421:23]
  wire [86:0] EmbeddedTLB_io_out_req_bits_user; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_out_resp_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_out_resp_valid; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 421:23]
  wire [86:0] EmbeddedTLB_io_out_resp_bits_user; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_mem_req_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 421:23]
  wire [31:0] EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 421:23]
  wire [3:0] EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_mem_resp_valid; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_flush; // @[EmbeddedTLB.scala 421:23]
  wire [1:0] EmbeddedTLB_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_cacheEmpty; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_io_ipf; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_CSRSATP; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_MOUFlushTLB; // @[EmbeddedTLB.scala 421:23]
  wire  Cache_clock; // @[Cache.scala 670:35]
  wire  Cache_reset; // @[Cache.scala 670:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 670:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 670:35]
  wire [86:0] Cache_io_in_req_bits_user; // @[Cache.scala 670:35]
  wire  Cache_io_in_resp_ready; // @[Cache.scala 670:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 670:35]
  wire [86:0] Cache_io_in_resp_bits_user; // @[Cache.scala 670:35]
  wire [1:0] Cache_io_flush; // @[Cache.scala 670:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 670:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 670:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 670:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 670:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 670:35]
  wire  Cache_io_mmio_req_ready; // @[Cache.scala 670:35]
  wire  Cache_io_mmio_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_io_mmio_req_bits_addr; // @[Cache.scala 670:35]
  wire  Cache_io_mmio_resp_valid; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_mmio_resp_bits_rdata; // @[Cache.scala 670:35]
  wire  Cache_io_empty; // @[Cache.scala 670:35]
  wire  Cache_MOUFlushICache; // @[Cache.scala 670:35]
  wire  EmbeddedTLB_1_clock; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_reset; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_in_req_valid; // @[EmbeddedTLB.scala 421:23]
  wire [38:0] EmbeddedTLB_1_io_in_req_bits_addr; // @[EmbeddedTLB.scala 421:23]
  wire [2:0] EmbeddedTLB_1_io_in_req_bits_size; // @[EmbeddedTLB.scala 421:23]
  wire [3:0] EmbeddedTLB_1_io_in_req_bits_cmd; // @[EmbeddedTLB.scala 421:23]
  wire [7:0] EmbeddedTLB_1_io_in_req_bits_wmask; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_1_io_in_req_bits_wdata; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_out_req_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_out_req_valid; // @[EmbeddedTLB.scala 421:23]
  wire [31:0] EmbeddedTLB_1_io_out_req_bits_addr; // @[EmbeddedTLB.scala 421:23]
  wire [2:0] EmbeddedTLB_1_io_out_req_bits_size; // @[EmbeddedTLB.scala 421:23]
  wire [3:0] EmbeddedTLB_1_io_out_req_bits_cmd; // @[EmbeddedTLB.scala 421:23]
  wire [7:0] EmbeddedTLB_1_io_out_req_bits_wmask; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_1_io_out_req_bits_wdata; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_out_resp_valid; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_1_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_mem_req_ready; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 421:23]
  wire [31:0] EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 421:23]
  wire [3:0] EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_mem_resp_valid; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_1_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 421:23]
  wire [1:0] EmbeddedTLB_1_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_sum; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 421:23]
  wire [38:0] EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1__T_28_0; // @[EmbeddedTLB.scala 421:23]
  wire [63:0] EmbeddedTLB_1_CSRSATP; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_amoReq; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_vmEnable_0; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1__T_27_0; // @[EmbeddedTLB.scala 421:23]
  wire  EmbeddedTLB_1_MOUFlushTLB; // @[EmbeddedTLB.scala 421:23]
  wire  Cache_1_clock; // @[Cache.scala 670:35]
  wire  Cache_1_reset; // @[Cache.scala 670:35]
  wire  Cache_1_io_in_req_ready; // @[Cache.scala 670:35]
  wire  Cache_1_io_in_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_1_io_in_req_bits_addr; // @[Cache.scala 670:35]
  wire [2:0] Cache_1_io_in_req_bits_size; // @[Cache.scala 670:35]
  wire [3:0] Cache_1_io_in_req_bits_cmd; // @[Cache.scala 670:35]
  wire [7:0] Cache_1_io_in_req_bits_wmask; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_in_req_bits_wdata; // @[Cache.scala 670:35]
  wire  Cache_1_io_in_resp_ready; // @[Cache.scala 670:35]
  wire  Cache_1_io_in_resp_valid; // @[Cache.scala 670:35]
  wire [3:0] Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 670:35]
  wire  Cache_1_io_out_mem_req_ready; // @[Cache.scala 670:35]
  wire  Cache_1_io_out_mem_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_1_io_out_mem_req_bits_addr; // @[Cache.scala 670:35]
  wire [3:0] Cache_1_io_out_mem_req_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_out_mem_req_bits_wdata; // @[Cache.scala 670:35]
  wire  Cache_1_io_out_mem_resp_valid; // @[Cache.scala 670:35]
  wire [3:0] Cache_1_io_out_mem_resp_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_out_mem_resp_bits_rdata; // @[Cache.scala 670:35]
  wire  Cache_1_io_out_coh_req_ready; // @[Cache.scala 670:35]
  wire  Cache_1_io_out_coh_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_1_io_out_coh_req_bits_addr; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_out_coh_req_bits_wdata; // @[Cache.scala 670:35]
  wire  Cache_1_io_out_coh_resp_valid; // @[Cache.scala 670:35]
  wire [3:0] Cache_1_io_out_coh_resp_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_out_coh_resp_bits_rdata; // @[Cache.scala 670:35]
  wire  Cache_1_io_mmio_req_ready; // @[Cache.scala 670:35]
  wire  Cache_1_io_mmio_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 670:35]
  wire [2:0] Cache_1_io_mmio_req_bits_size; // @[Cache.scala 670:35]
  wire [3:0] Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 670:35]
  wire [7:0] Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 670:35]
  wire  Cache_1_io_mmio_resp_valid; // @[Cache.scala 670:35]
  wire [63:0] Cache_1_io_mmio_resp_bits_rdata; // @[Cache.scala 670:35]
  reg [63:0] REG__0_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__0_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__0_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__0_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__0_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__0_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__0_ctrl_vtag; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_vec_addr; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__0_ctrl_length_k; // @[PipelineVector.scala 29:29]
  reg [1:0] REG__0_ctrl_algorithm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__0_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__1_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__1_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__1_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__1_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__1_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__1_ctrl_vtag; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_vec_addr; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__1_ctrl_length_k; // @[PipelineVector.scala 29:29]
  reg [1:0] REG__1_ctrl_algorithm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__2_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__2_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__2_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__2_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__2_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__2_ctrl_vtag; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_vec_addr; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__2_ctrl_length_k; // @[PipelineVector.scala 29:29]
  reg [1:0] REG__2_ctrl_algorithm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__3_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__3_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__3_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__3_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__3_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__3_ctrl_vtag; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_vec_addr; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__3_ctrl_length_k; // @[PipelineVector.scala 29:29]
  reg [1:0] REG__3_ctrl_algorithm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_data_imm; // @[PipelineVector.scala 29:29]
  reg [1:0] REG_1; // @[PipelineVector.scala 30:33]
  reg [1:0] REG_2; // @[PipelineVector.scala 31:33]
  wire [1:0] _T_3 = REG_1 + 2'h1; // @[PipelineVector.scala 33:63]
  wire [1:0] _T_6 = REG_1 + 2'h2; // @[PipelineVector.scala 33:63]
  wire  _T_9 = _T_3 != REG_2 & _T_6 != REG_2; // @[PipelineVector.scala 33:124]
  wire  _WIRE_5_0 = frontend_io_out_0_valid; // @[PipelineVector.scala 36:27 37:20]
  wire  _WIRE_5_1 = frontend_io_out_1_valid; // @[PipelineVector.scala 36:27 38:20]
  wire [1:0] _T_10 = _WIRE_5_0 + _WIRE_5_1; // @[PipelineVector.scala 40:46]
  wire  _T_11 = _T_10 >= 2'h1; // @[PipelineVector.scala 41:53]
  wire  _T_12 = _T_10 >= 2'h2; // @[PipelineVector.scala 41:53]
  wire  _T_13 = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = frontend_io_out_1_ready & frontend_io_out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_15 = _T_13 | _T_14; // @[PipelineVector.scala 43:26]
  wire [2:0] _T_16 = {{1'd0}, REG_1}; // @[PipelineVector.scala 45:45]
  wire [63:0] _T_18_cf_instr = _WIRE_5_0 ? frontend_io_out_0_bits_cf_instr : frontend_io_out_1_bits_cf_instr; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_18_cf_pc = _WIRE_5_0 ? frontend_io_out_0_bits_cf_pc : frontend_io_out_1_bits_cf_pc; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_18_cf_pnpc = _WIRE_5_0 ? frontend_io_out_0_bits_cf_pnpc : frontend_io_out_1_bits_cf_pnpc; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_exceptionVec_1 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_exceptionVec_1 :
    frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_exceptionVec_2 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_exceptionVec_2 :
    frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_exceptionVec_12 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_exceptionVec_12 :
    frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_0 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_0 : frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_1 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_1 : frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_2 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_2 : frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_3 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_3 : frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_4 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_4 : frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_5 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_5 : frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_6 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_6 : frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_7 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_7 : frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_8 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_8 : frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_9 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_9 : frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_10 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_10 : frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_11 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_11 : frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 45:69]
  wire [3:0] _T_18_cf_brIdx = _WIRE_5_0 ? frontend_io_out_0_bits_cf_brIdx : frontend_io_out_1_bits_cf_brIdx; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_crossPageIPFFix = _WIRE_5_0 ? frontend_io_out_0_bits_cf_crossPageIPFFix :
    frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 45:69]
  wire [63:0] _T_18_cf_runahead_checkpoint_id = _WIRE_5_0 ? frontend_io_out_0_bits_cf_runahead_checkpoint_id : 64'h0; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_src1Type = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_src1Type : frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_src2Type = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_src2Type : frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 45:69]
  wire [2:0] _T_18_ctrl_fuType = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_fuType : frontend_io_out_1_bits_ctrl_fuType; // @[PipelineVector.scala 45:69]
  wire [6:0] _T_18_ctrl_fuOpType = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_fuOpType :
    frontend_io_out_1_bits_ctrl_fuOpType; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfSrc1 = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : frontend_io_out_1_bits_ctrl_rfSrc1; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfSrc2 = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : frontend_io_out_1_bits_ctrl_rfSrc2; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_rfWen = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfWen : frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfDest = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfDest : frontend_io_out_1_bits_ctrl_rfDest; // @[PipelineVector.scala 45:69]
  wire [2:0] _T_18_ctrl_vtag = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_vtag : frontend_io_out_1_bits_ctrl_vtag; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_vec_addr = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_vec_addr :
    frontend_io_out_1_bits_ctrl_vec_addr; // @[PipelineVector.scala 45:69]
  wire [3:0] _T_18_ctrl_length_k = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_length_k :
    frontend_io_out_1_bits_ctrl_length_k; // @[PipelineVector.scala 45:69]
  wire [1:0] _T_18_ctrl_algorithm = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_algorithm :
    frontend_io_out_1_bits_ctrl_algorithm; // @[PipelineVector.scala 45:69]
  wire [63:0] _T_18_data_imm = _WIRE_5_0 ? frontend_io_out_0_bits_data_imm : frontend_io_out_1_bits_data_imm; // @[PipelineVector.scala 45:69]
  wire [63:0] _GEN_0 = 2'h0 == _T_16[1:0] ? _T_18_data_imm : REG__0_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_1 = 2'h1 == _T_16[1:0] ? _T_18_data_imm : REG__1_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_2 = 2'h2 == _T_16[1:0] ? _T_18_data_imm : REG__2_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_3 = 2'h3 == _T_16[1:0] ? _T_18_data_imm : REG__3_data_imm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [1:0] _GEN_12 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_algorithm : REG__0_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [1:0] _GEN_13 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_algorithm : REG__1_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [1:0] _GEN_14 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_algorithm : REG__2_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [1:0] _GEN_15 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_algorithm : REG__3_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_16 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_length_k : REG__0_ctrl_length_k; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_17 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_length_k : REG__1_ctrl_length_k; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_18 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_length_k : REG__2_ctrl_length_k; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_19 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_length_k : REG__3_ctrl_length_k; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_20 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_vec_addr : REG__0_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_21 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_vec_addr : REG__1_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_22 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_vec_addr : REG__2_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_23 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_vec_addr : REG__3_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_24 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_vtag : REG__0_ctrl_vtag; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_25 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_vtag : REG__1_ctrl_vtag; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_26 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_vtag : REG__2_ctrl_vtag; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_27 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_vtag : REG__3_ctrl_vtag; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_48 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__0_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_49 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__1_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_50 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__2_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_51 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__3_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_52 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__0_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_53 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__1_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_54 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__2_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_55 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__3_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_56 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_57 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_58 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_59 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_60 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_61 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_62 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_63 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_64 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_65 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__1_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_66 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__2_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_67 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__3_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_68 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__0_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_69 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__1_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_70 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__2_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_71 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__3_ctrl_fuType; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_72 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__0_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_73 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__1_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_74 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__2_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_75 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__3_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_76 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__0_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_77 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__1_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_78 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__2_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_79 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__3_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_84 = 2'h0 == _T_16[1:0] ? _T_18_cf_runahead_checkpoint_id : REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_85 = 2'h1 == _T_16[1:0] ? _T_18_cf_runahead_checkpoint_id : REG__1_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_86 = 2'h2 == _T_16[1:0] ? _T_18_cf_runahead_checkpoint_id : REG__2_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_87 = 2'h3 == _T_16[1:0] ? _T_18_cf_runahead_checkpoint_id : REG__3_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_88 = 2'h0 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_89 = 2'h1 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_90 = 2'h2 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_91 = 2'h3 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_96 = 2'h0 == _T_16[1:0] ? _T_18_cf_brIdx : REG__0_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_97 = 2'h1 == _T_16[1:0] ? _T_18_cf_brIdx : REG__1_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_98 = 2'h2 == _T_16[1:0] ? _T_18_cf_brIdx : REG__2_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_99 = 2'h3 == _T_16[1:0] ? _T_18_cf_brIdx : REG__3_cf_brIdx; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_100 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_101 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__1_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_102 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__2_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_103 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__3_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_104 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_105 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__1_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_106 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__2_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_107 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__3_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_108 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_109 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__1_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_110 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__2_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_111 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__3_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_112 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_113 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__1_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_114 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__2_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_115 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__3_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_116 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_117 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__1_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_118 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__2_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_119 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__3_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_120 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_121 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__1_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_122 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__2_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_123 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__3_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_124 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_125 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__1_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_126 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__2_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_127 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__3_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_128 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_129 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__1_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_130 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__2_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_131 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__3_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_132 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_133 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__1_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_134 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__2_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_135 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__3_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_136 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_137 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__1_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_138 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__2_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_139 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__3_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_140 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_141 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__1_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_142 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__2_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_143 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__3_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_144 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_145 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__1_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_146 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__2_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_147 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__3_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_152 = 2'h0 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_153 = 2'h1 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_154 = 2'h2 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_155 = 2'h3 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_156 = 2'h0 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_157 = 2'h1 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_158 = 2'h2 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_159 = 2'h3 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_196 = 2'h0 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_197 = 2'h1 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_198 = 2'h2 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_199 = 2'h3 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_224 = 2'h0 == _T_16[1:0] ? _T_18_cf_pnpc : REG__0_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_225 = 2'h1 == _T_16[1:0] ? _T_18_cf_pnpc : REG__1_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_226 = 2'h2 == _T_16[1:0] ? _T_18_cf_pnpc : REG__2_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_227 = 2'h3 == _T_16[1:0] ? _T_18_cf_pnpc : REG__3_cf_pnpc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_228 = 2'h0 == _T_16[1:0] ? _T_18_cf_pc : REG__0_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_229 = 2'h1 == _T_16[1:0] ? _T_18_cf_pc : REG__1_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_230 = 2'h2 == _T_16[1:0] ? _T_18_cf_pc : REG__2_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_231 = 2'h3 == _T_16[1:0] ? _T_18_cf_pc : REG__3_cf_pc; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_232 = 2'h0 == _T_16[1:0] ? _T_18_cf_instr : REG__0_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_233 = 2'h1 == _T_16[1:0] ? _T_18_cf_instr : REG__1_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_234 = 2'h2 == _T_16[1:0] ? _T_18_cf_instr : REG__2_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_235 = 2'h3 == _T_16[1:0] ? _T_18_cf_instr : REG__3_cf_instr; // @[PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_236 = _T_11 ? _GEN_0 : REG__0_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_237 = _T_11 ? _GEN_1 : REG__1_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_238 = _T_11 ? _GEN_2 : REG__2_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_239 = _T_11 ? _GEN_3 : REG__3_data_imm; // @[PipelineVector.scala 29:29 45:29]
  wire [1:0] _GEN_248 = _T_11 ? _GEN_12 : REG__0_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:29]
  wire [1:0] _GEN_249 = _T_11 ? _GEN_13 : REG__1_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:29]
  wire [1:0] _GEN_250 = _T_11 ? _GEN_14 : REG__2_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:29]
  wire [1:0] _GEN_251 = _T_11 ? _GEN_15 : REG__3_ctrl_algorithm; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_252 = _T_11 ? _GEN_16 : REG__0_ctrl_length_k; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_253 = _T_11 ? _GEN_17 : REG__1_ctrl_length_k; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_254 = _T_11 ? _GEN_18 : REG__2_ctrl_length_k; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_255 = _T_11 ? _GEN_19 : REG__3_ctrl_length_k; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_256 = _T_11 ? _GEN_20 : REG__0_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_257 = _T_11 ? _GEN_21 : REG__1_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_258 = _T_11 ? _GEN_22 : REG__2_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_259 = _T_11 ? _GEN_23 : REG__3_ctrl_vec_addr; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_260 = _T_11 ? _GEN_24 : REG__0_ctrl_vtag; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_261 = _T_11 ? _GEN_25 : REG__1_ctrl_vtag; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_262 = _T_11 ? _GEN_26 : REG__2_ctrl_vtag; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_263 = _T_11 ? _GEN_27 : REG__3_ctrl_vtag; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_284 = _T_11 ? _GEN_48 : REG__0_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_285 = _T_11 ? _GEN_49 : REG__1_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_286 = _T_11 ? _GEN_50 : REG__2_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_287 = _T_11 ? _GEN_51 : REG__3_ctrl_rfDest; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_288 = _T_11 ? _GEN_52 : REG__0_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_289 = _T_11 ? _GEN_53 : REG__1_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_290 = _T_11 ? _GEN_54 : REG__2_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_291 = _T_11 ? _GEN_55 : REG__3_ctrl_rfWen; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_292 = _T_11 ? _GEN_56 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_293 = _T_11 ? _GEN_57 : REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_294 = _T_11 ? _GEN_58 : REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_295 = _T_11 ? _GEN_59 : REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_296 = _T_11 ? _GEN_60 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_297 = _T_11 ? _GEN_61 : REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_298 = _T_11 ? _GEN_62 : REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_299 = _T_11 ? _GEN_63 : REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_300 = _T_11 ? _GEN_64 : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_301 = _T_11 ? _GEN_65 : REG__1_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_302 = _T_11 ? _GEN_66 : REG__2_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_303 = _T_11 ? _GEN_67 : REG__3_ctrl_fuOpType; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_304 = _T_11 ? _GEN_68 : REG__0_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_305 = _T_11 ? _GEN_69 : REG__1_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_306 = _T_11 ? _GEN_70 : REG__2_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_307 = _T_11 ? _GEN_71 : REG__3_ctrl_fuType; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_308 = _T_11 ? _GEN_72 : REG__0_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_309 = _T_11 ? _GEN_73 : REG__1_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_310 = _T_11 ? _GEN_74 : REG__2_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_311 = _T_11 ? _GEN_75 : REG__3_ctrl_src2Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_312 = _T_11 ? _GEN_76 : REG__0_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_313 = _T_11 ? _GEN_77 : REG__1_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_314 = _T_11 ? _GEN_78 : REG__2_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_315 = _T_11 ? _GEN_79 : REG__3_ctrl_src1Type; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_320 = _T_11 ? _GEN_84 : REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_321 = _T_11 ? _GEN_85 : REG__1_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_322 = _T_11 ? _GEN_86 : REG__2_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_323 = _T_11 ? _GEN_87 : REG__3_cf_runahead_checkpoint_id; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_324 = _T_11 ? _GEN_88 : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_325 = _T_11 ? _GEN_89 : REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_326 = _T_11 ? _GEN_90 : REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_327 = _T_11 ? _GEN_91 : REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_332 = _T_11 ? _GEN_96 : REG__0_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_333 = _T_11 ? _GEN_97 : REG__1_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_334 = _T_11 ? _GEN_98 : REG__2_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_335 = _T_11 ? _GEN_99 : REG__3_cf_brIdx; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_336 = _T_11 ? _GEN_100 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_337 = _T_11 ? _GEN_101 : REG__1_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_338 = _T_11 ? _GEN_102 : REG__2_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_339 = _T_11 ? _GEN_103 : REG__3_cf_intrVec_0; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_340 = _T_11 ? _GEN_104 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_341 = _T_11 ? _GEN_105 : REG__1_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_342 = _T_11 ? _GEN_106 : REG__2_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_343 = _T_11 ? _GEN_107 : REG__3_cf_intrVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_344 = _T_11 ? _GEN_108 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_345 = _T_11 ? _GEN_109 : REG__1_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_346 = _T_11 ? _GEN_110 : REG__2_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_347 = _T_11 ? _GEN_111 : REG__3_cf_intrVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_348 = _T_11 ? _GEN_112 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_349 = _T_11 ? _GEN_113 : REG__1_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_350 = _T_11 ? _GEN_114 : REG__2_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_351 = _T_11 ? _GEN_115 : REG__3_cf_intrVec_3; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_352 = _T_11 ? _GEN_116 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_353 = _T_11 ? _GEN_117 : REG__1_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_354 = _T_11 ? _GEN_118 : REG__2_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_355 = _T_11 ? _GEN_119 : REG__3_cf_intrVec_4; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_356 = _T_11 ? _GEN_120 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_357 = _T_11 ? _GEN_121 : REG__1_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_358 = _T_11 ? _GEN_122 : REG__2_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_359 = _T_11 ? _GEN_123 : REG__3_cf_intrVec_5; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_360 = _T_11 ? _GEN_124 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_361 = _T_11 ? _GEN_125 : REG__1_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_362 = _T_11 ? _GEN_126 : REG__2_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_363 = _T_11 ? _GEN_127 : REG__3_cf_intrVec_6; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_364 = _T_11 ? _GEN_128 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_365 = _T_11 ? _GEN_129 : REG__1_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_366 = _T_11 ? _GEN_130 : REG__2_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_367 = _T_11 ? _GEN_131 : REG__3_cf_intrVec_7; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_368 = _T_11 ? _GEN_132 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_369 = _T_11 ? _GEN_133 : REG__1_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_370 = _T_11 ? _GEN_134 : REG__2_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_371 = _T_11 ? _GEN_135 : REG__3_cf_intrVec_8; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_372 = _T_11 ? _GEN_136 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_373 = _T_11 ? _GEN_137 : REG__1_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_374 = _T_11 ? _GEN_138 : REG__2_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_375 = _T_11 ? _GEN_139 : REG__3_cf_intrVec_9; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_376 = _T_11 ? _GEN_140 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_377 = _T_11 ? _GEN_141 : REG__1_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_378 = _T_11 ? _GEN_142 : REG__2_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_379 = _T_11 ? _GEN_143 : REG__3_cf_intrVec_10; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_380 = _T_11 ? _GEN_144 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_381 = _T_11 ? _GEN_145 : REG__1_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_382 = _T_11 ? _GEN_146 : REG__2_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_383 = _T_11 ? _GEN_147 : REG__3_cf_intrVec_11; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_388 = _T_11 ? _GEN_152 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_389 = _T_11 ? _GEN_153 : REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_390 = _T_11 ? _GEN_154 : REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_391 = _T_11 ? _GEN_155 : REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_392 = _T_11 ? _GEN_156 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_393 = _T_11 ? _GEN_157 : REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_394 = _T_11 ? _GEN_158 : REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_395 = _T_11 ? _GEN_159 : REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_432 = _T_11 ? _GEN_196 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_433 = _T_11 ? _GEN_197 : REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_434 = _T_11 ? _GEN_198 : REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire  _GEN_435 = _T_11 ? _GEN_199 : REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_460 = _T_11 ? _GEN_224 : REG__0_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_461 = _T_11 ? _GEN_225 : REG__1_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_462 = _T_11 ? _GEN_226 : REG__2_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_463 = _T_11 ? _GEN_227 : REG__3_cf_pnpc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_464 = _T_11 ? _GEN_228 : REG__0_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_465 = _T_11 ? _GEN_229 : REG__1_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_466 = _T_11 ? _GEN_230 : REG__2_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_467 = _T_11 ? _GEN_231 : REG__3_cf_pc; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_468 = _T_11 ? _GEN_232 : REG__0_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_469 = _T_11 ? _GEN_233 : REG__1_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_470 = _T_11 ? _GEN_234 : REG__2_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_471 = _T_11 ? _GEN_235 : REG__3_cf_instr; // @[PipelineVector.scala 29:29 45:29]
  wire [1:0] _T_20 = 2'h1 + REG_1; // @[PipelineVector.scala 46:45]
  wire [63:0] _REG_T_20_data_imm = frontend_io_out_1_bits_data_imm; // @[PipelineVector.scala 46:{63,63}]
  wire [1:0] _REG_T_20_ctrl_algorithm = frontend_io_out_1_bits_ctrl_algorithm; // @[PipelineVector.scala 46:{63,63}]
  wire [3:0] _REG_T_20_ctrl_length_k = frontend_io_out_1_bits_ctrl_length_k; // @[PipelineVector.scala 46:{63,63}]
  wire [4:0] _REG_T_20_ctrl_vec_addr = frontend_io_out_1_bits_ctrl_vec_addr; // @[PipelineVector.scala 46:{63,63}]
  wire [2:0] _REG_T_20_ctrl_vtag = frontend_io_out_1_bits_ctrl_vtag; // @[PipelineVector.scala 46:{63,63}]
  wire [4:0] _REG_T_20_ctrl_rfDest = frontend_io_out_1_bits_ctrl_rfDest; // @[PipelineVector.scala 46:{63,63}]
  wire [4:0] _REG_T_20_ctrl_rfSrc2 = frontend_io_out_1_bits_ctrl_rfSrc2; // @[PipelineVector.scala 46:{63,63}]
  wire [4:0] _REG_T_20_ctrl_rfSrc1 = frontend_io_out_1_bits_ctrl_rfSrc1; // @[PipelineVector.scala 46:{63,63}]
  wire [6:0] _REG_T_20_ctrl_fuOpType = frontend_io_out_1_bits_ctrl_fuOpType; // @[PipelineVector.scala 46:{63,63}]
  wire [2:0] _REG_T_20_ctrl_fuType = frontend_io_out_1_bits_ctrl_fuType; // @[PipelineVector.scala 46:{63,63}]
  wire [3:0] _REG_T_20_cf_brIdx = frontend_io_out_1_bits_cf_brIdx; // @[PipelineVector.scala 46:{63,63}]
  wire [38:0] _REG_T_20_cf_pnpc = frontend_io_out_1_bits_cf_pnpc; // @[PipelineVector.scala 46:{63,63}]
  wire [38:0] _REG_T_20_cf_pc = frontend_io_out_1_bits_cf_pc; // @[PipelineVector.scala 46:{63,63}]
  wire [63:0] _REG_T_20_cf_instr = frontend_io_out_1_bits_cf_instr; // @[PipelineVector.scala 46:{63,63}]
  wire [1:0] _T_22 = REG_1 + _T_10; // @[PipelineVector.scala 47:42]
  wire [63:0] _GEN_1182 = 2'h1 == REG_2 ? REG__1_data_imm : REG__0_data_imm; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1183 = 2'h2 == REG_2 ? REG__2_data_imm : _GEN_1182; // @[PipelineVector.scala 55:{15,15}]
  wire [1:0] _GEN_1194 = 2'h1 == REG_2 ? REG__1_ctrl_algorithm : REG__0_ctrl_algorithm; // @[PipelineVector.scala 55:{15,15}]
  wire [1:0] _GEN_1195 = 2'h2 == REG_2 ? REG__2_ctrl_algorithm : _GEN_1194; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1198 = 2'h1 == REG_2 ? REG__1_ctrl_length_k : REG__0_ctrl_length_k; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1199 = 2'h2 == REG_2 ? REG__2_ctrl_length_k : _GEN_1198; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1202 = 2'h1 == REG_2 ? REG__1_ctrl_vec_addr : REG__0_ctrl_vec_addr; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1203 = 2'h2 == REG_2 ? REG__2_ctrl_vec_addr : _GEN_1202; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1206 = 2'h1 == REG_2 ? REG__1_ctrl_vtag : REG__0_ctrl_vtag; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1207 = 2'h2 == REG_2 ? REG__2_ctrl_vtag : _GEN_1206; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1230 = 2'h1 == REG_2 ? REG__1_ctrl_rfDest : REG__0_ctrl_rfDest; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1231 = 2'h2 == REG_2 ? REG__2_ctrl_rfDest : _GEN_1230; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1234 = 2'h1 == REG_2 ? REG__1_ctrl_rfWen : REG__0_ctrl_rfWen; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1235 = 2'h2 == REG_2 ? REG__2_ctrl_rfWen : _GEN_1234; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1238 = 2'h1 == REG_2 ? REG__1_ctrl_rfSrc2 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1239 = 2'h2 == REG_2 ? REG__2_ctrl_rfSrc2 : _GEN_1238; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1242 = 2'h1 == REG_2 ? REG__1_ctrl_rfSrc1 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1243 = 2'h2 == REG_2 ? REG__2_ctrl_rfSrc1 : _GEN_1242; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1246 = 2'h1 == REG_2 ? REG__1_ctrl_fuOpType : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1247 = 2'h2 == REG_2 ? REG__2_ctrl_fuOpType : _GEN_1246; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1250 = 2'h1 == REG_2 ? REG__1_ctrl_fuType : REG__0_ctrl_fuType; // @[PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1251 = 2'h2 == REG_2 ? REG__2_ctrl_fuType : _GEN_1250; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1254 = 2'h1 == REG_2 ? REG__1_ctrl_src2Type : REG__0_ctrl_src2Type; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1255 = 2'h2 == REG_2 ? REG__2_ctrl_src2Type : _GEN_1254; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1258 = 2'h1 == REG_2 ? REG__1_ctrl_src1Type : REG__0_ctrl_src1Type; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1259 = 2'h2 == REG_2 ? REG__2_ctrl_src1Type : _GEN_1258; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1266 = 2'h1 == REG_2 ? REG__1_cf_runahead_checkpoint_id : REG__0_cf_runahead_checkpoint_id; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1267 = 2'h2 == REG_2 ? REG__2_cf_runahead_checkpoint_id : _GEN_1266; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1270 = 2'h1 == REG_2 ? REG__1_cf_crossPageIPFFix : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1271 = 2'h2 == REG_2 ? REG__2_cf_crossPageIPFFix : _GEN_1270; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1278 = 2'h1 == REG_2 ? REG__1_cf_brIdx : REG__0_cf_brIdx; // @[PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1279 = 2'h2 == REG_2 ? REG__2_cf_brIdx : _GEN_1278; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1282 = 2'h1 == REG_2 ? REG__1_cf_intrVec_0 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1283 = 2'h2 == REG_2 ? REG__2_cf_intrVec_0 : _GEN_1282; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1286 = 2'h1 == REG_2 ? REG__1_cf_intrVec_1 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1287 = 2'h2 == REG_2 ? REG__2_cf_intrVec_1 : _GEN_1286; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1290 = 2'h1 == REG_2 ? REG__1_cf_intrVec_2 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1291 = 2'h2 == REG_2 ? REG__2_cf_intrVec_2 : _GEN_1290; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1294 = 2'h1 == REG_2 ? REG__1_cf_intrVec_3 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1295 = 2'h2 == REG_2 ? REG__2_cf_intrVec_3 : _GEN_1294; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1298 = 2'h1 == REG_2 ? REG__1_cf_intrVec_4 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1299 = 2'h2 == REG_2 ? REG__2_cf_intrVec_4 : _GEN_1298; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1302 = 2'h1 == REG_2 ? REG__1_cf_intrVec_5 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1303 = 2'h2 == REG_2 ? REG__2_cf_intrVec_5 : _GEN_1302; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1306 = 2'h1 == REG_2 ? REG__1_cf_intrVec_6 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1307 = 2'h2 == REG_2 ? REG__2_cf_intrVec_6 : _GEN_1306; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1310 = 2'h1 == REG_2 ? REG__1_cf_intrVec_7 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1311 = 2'h2 == REG_2 ? REG__2_cf_intrVec_7 : _GEN_1310; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1314 = 2'h1 == REG_2 ? REG__1_cf_intrVec_8 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1315 = 2'h2 == REG_2 ? REG__2_cf_intrVec_8 : _GEN_1314; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1318 = 2'h1 == REG_2 ? REG__1_cf_intrVec_9 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1319 = 2'h2 == REG_2 ? REG__2_cf_intrVec_9 : _GEN_1318; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1322 = 2'h1 == REG_2 ? REG__1_cf_intrVec_10 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1323 = 2'h2 == REG_2 ? REG__2_cf_intrVec_10 : _GEN_1322; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1326 = 2'h1 == REG_2 ? REG__1_cf_intrVec_11 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1327 = 2'h2 == REG_2 ? REG__2_cf_intrVec_11 : _GEN_1326; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1334 = 2'h1 == REG_2 ? REG__1_cf_exceptionVec_1 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1335 = 2'h2 == REG_2 ? REG__2_cf_exceptionVec_1 : _GEN_1334; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1338 = 2'h1 == REG_2 ? REG__1_cf_exceptionVec_2 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1339 = 2'h2 == REG_2 ? REG__2_cf_exceptionVec_2 : _GEN_1338; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1378 = 2'h1 == REG_2 ? REG__1_cf_exceptionVec_12 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 55:{15,15}]
  wire  _GEN_1379 = 2'h2 == REG_2 ? REG__2_cf_exceptionVec_12 : _GEN_1378; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1406 = 2'h1 == REG_2 ? REG__1_cf_pnpc : REG__0_cf_pnpc; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1407 = 2'h2 == REG_2 ? REG__2_cf_pnpc : _GEN_1406; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1410 = 2'h1 == REG_2 ? REG__1_cf_pc : REG__0_cf_pc; // @[PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1411 = 2'h2 == REG_2 ? REG__2_cf_pc : _GEN_1410; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1414 = 2'h1 == REG_2 ? REG__1_cf_instr : REG__0_cf_instr; // @[PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1415 = 2'h2 == REG_2 ? REG__2_cf_instr : _GEN_1414; // @[PipelineVector.scala 55:{15,15}]
  wire  _T_32 = Backend_inorder_io_in_0_ready & Backend_inorder_io_in_0_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_34 = {{1'd0}, _T_32}; // @[PipelineVector.scala 64:44]
  wire  _T_35 = _T_34 > 2'h0; // @[PipelineVector.scala 65:35]
  wire [1:0] _T_37 = REG_2 + _T_34; // @[PipelineVector.scala 67:42]
  Frontend_inorder frontend ( // @[NutCore.scala 104:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(frontend_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(frontend_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(frontend_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(frontend_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(frontend_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(frontend_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(frontend_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_cf_runahead_checkpoint_id(frontend_io_out_0_bits_cf_runahead_checkpoint_id),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_vtag(frontend_io_out_0_bits_ctrl_vtag),
    .io_out_0_bits_ctrl_vec_addr(frontend_io_out_0_bits_ctrl_vec_addr),
    .io_out_0_bits_ctrl_length_k(frontend_io_out_0_bits_ctrl_length_k),
    .io_out_0_bits_ctrl_algorithm(frontend_io_out_0_bits_ctrl_algorithm),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_out_1_ready(frontend_io_out_1_ready),
    .io_out_1_valid(frontend_io_out_1_valid),
    .io_out_1_bits_cf_instr(frontend_io_out_1_bits_cf_instr),
    .io_out_1_bits_cf_pc(frontend_io_out_1_bits_cf_pc),
    .io_out_1_bits_cf_pnpc(frontend_io_out_1_bits_cf_pnpc),
    .io_out_1_bits_cf_exceptionVec_1(frontend_io_out_1_bits_cf_exceptionVec_1),
    .io_out_1_bits_cf_exceptionVec_2(frontend_io_out_1_bits_cf_exceptionVec_2),
    .io_out_1_bits_cf_exceptionVec_12(frontend_io_out_1_bits_cf_exceptionVec_12),
    .io_out_1_bits_cf_intrVec_0(frontend_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(frontend_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(frontend_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(frontend_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(frontend_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(frontend_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(frontend_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(frontend_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(frontend_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(frontend_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(frontend_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(frontend_io_out_1_bits_cf_intrVec_11),
    .io_out_1_bits_cf_brIdx(frontend_io_out_1_bits_cf_brIdx),
    .io_out_1_bits_cf_crossPageIPFFix(frontend_io_out_1_bits_cf_crossPageIPFFix),
    .io_out_1_bits_ctrl_src1Type(frontend_io_out_1_bits_ctrl_src1Type),
    .io_out_1_bits_ctrl_src2Type(frontend_io_out_1_bits_ctrl_src2Type),
    .io_out_1_bits_ctrl_fuType(frontend_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(frontend_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_rfSrc1(frontend_io_out_1_bits_ctrl_rfSrc1),
    .io_out_1_bits_ctrl_rfSrc2(frontend_io_out_1_bits_ctrl_rfSrc2),
    .io_out_1_bits_ctrl_rfWen(frontend_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_rfDest(frontend_io_out_1_bits_ctrl_rfDest),
    .io_out_1_bits_ctrl_vtag(frontend_io_out_1_bits_ctrl_vtag),
    .io_out_1_bits_ctrl_vec_addr(frontend_io_out_1_bits_ctrl_vec_addr),
    .io_out_1_bits_ctrl_length_k(frontend_io_out_1_bits_ctrl_length_k),
    .io_out_1_bits_ctrl_algorithm(frontend_io_out_1_bits_ctrl_algorithm),
    .io_out_1_bits_data_imm(frontend_io_out_1_bits_data_imm),
    .io_flushVec(frontend_io_flushVec),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .io_ipf(frontend_io_ipf),
    .flushICache(frontend_flushICache),
    .REG_0_valid(frontend_REG_0_valid),
    .REG_0_pc(frontend_REG_0_pc),
    .REG_0_isMissPredict(frontend_REG_0_isMissPredict),
    .REG_0_actualTarget(frontend_REG_0_actualTarget),
    .REG_0_actualTaken(frontend_REG_0_actualTaken),
    .REG_0_fuOpType(frontend_REG_0_fuOpType),
    .REG_0_btbType(frontend_REG_0_btbType),
    .REG_0_isRVC(frontend_REG_0_isRVC),
    .vmEnable(frontend_vmEnable),
    .intrVec(frontend_intrVec),
    .flushTLB(frontend_flushTLB)
  );
  Backend_inorder Backend_inorder ( // @[NutCore.scala 147:25]
    .clock(Backend_inorder_clock),
    .reset(Backend_inorder_reset),
    .io_in_0_ready(Backend_inorder_io_in_0_ready),
    .io_in_0_valid(Backend_inorder_io_in_0_valid),
    .io_in_0_bits_cf_instr(Backend_inorder_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(Backend_inorder_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(Backend_inorder_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(Backend_inorder_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(Backend_inorder_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(Backend_inorder_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(Backend_inorder_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(Backend_inorder_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(Backend_inorder_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(Backend_inorder_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(Backend_inorder_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(Backend_inorder_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(Backend_inorder_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(Backend_inorder_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(Backend_inorder_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(Backend_inorder_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(Backend_inorder_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(Backend_inorder_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(Backend_inorder_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(Backend_inorder_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_cf_runahead_checkpoint_id(Backend_inorder_io_in_0_bits_cf_runahead_checkpoint_id),
    .io_in_0_bits_ctrl_src1Type(Backend_inorder_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(Backend_inorder_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(Backend_inorder_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(Backend_inorder_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(Backend_inorder_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(Backend_inorder_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(Backend_inorder_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(Backend_inorder_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_vtag(Backend_inorder_io_in_0_bits_ctrl_vtag),
    .io_in_0_bits_ctrl_vec_addr(Backend_inorder_io_in_0_bits_ctrl_vec_addr),
    .io_in_0_bits_ctrl_length_k(Backend_inorder_io_in_0_bits_ctrl_length_k),
    .io_in_0_bits_ctrl_algorithm(Backend_inorder_io_in_0_bits_ctrl_algorithm),
    .io_in_0_bits_data_imm(Backend_inorder_io_in_0_bits_data_imm),
    .io_flush(Backend_inorder_io_flush),
    .io_dmem_req_ready(Backend_inorder_io_dmem_req_ready),
    .io_dmem_req_valid(Backend_inorder_io_dmem_req_valid),
    .io_dmem_req_bits_addr(Backend_inorder_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(Backend_inorder_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(Backend_inorder_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(Backend_inorder_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(Backend_inorder_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(Backend_inorder_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(Backend_inorder_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(Backend_inorder_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(Backend_inorder_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(Backend_inorder_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(Backend_inorder_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(Backend_inorder_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(Backend_inorder_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_addr(Backend_inorder_io_memMMU_dmem_addr),
    .io_redirect_target(Backend_inorder_io_redirect_target),
    .io_redirect_valid(Backend_inorder_io_redirect_valid),
    ._T_28(Backend_inorder__T_28),
    .flushICache(Backend_inorder_flushICache),
    .perfCnts_2(Backend_inorder_perfCnts_2),
    .io_in_bits_decode_cf_pc(Backend_inorder_io_in_bits_decode_cf_pc),
    .satp(Backend_inorder_satp),
    .REG_0_valid(Backend_inorder_REG_0_valid),
    .REG_0_pc(Backend_inorder_REG_0_pc),
    .REG_0_isMissPredict(Backend_inorder_REG_0_isMissPredict),
    .REG_0_actualTarget(Backend_inorder_REG_0_actualTarget),
    .REG_0_actualTaken(Backend_inorder_REG_0_actualTaken),
    .REG_0_fuOpType(Backend_inorder_REG_0_fuOpType),
    .REG_0_btbType(Backend_inorder_REG_0_btbType),
    .REG_0_isRVC(Backend_inorder_REG_0_isRVC),
    .io_wb_rfDest(Backend_inorder_io_wb_rfDest),
    .io_extra_mtip(Backend_inorder_io_extra_mtip),
    .amoReq(Backend_inorder_amoReq),
    .io_extra_meip_0(Backend_inorder_io_extra_meip_0),
    .vmEnable(Backend_inorder_vmEnable),
    .io_wb_rfWen(Backend_inorder_io_wb_rfWen),
    .io_wb_rfData(Backend_inorder_io_wb_rfData),
    .intrVec(Backend_inorder_intrVec),
    ._T_27(Backend_inorder__T_27),
    .io_extra_msip(Backend_inorder_io_extra_msip),
    .flushTLB(Backend_inorder_flushTLB),
    .io_in_valid_0(Backend_inorder_io_in_valid_0)
  );
  SimpleBusCrossbarNto1 SimpleBusCrossbarNto1 ( // @[NutCore.scala 151:26]
    .clock(SimpleBusCrossbarNto1_clock),
    .reset(SimpleBusCrossbarNto1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(SimpleBusCrossbarNto1_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(SimpleBusCrossbarNto1_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 SimpleBusCrossbarNto1_1 ( // @[NutCore.scala 152:26]
    .clock(SimpleBusCrossbarNto1_1_clock),
    .reset(SimpleBusCrossbarNto1_1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(SimpleBusCrossbarNto1_1_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_1_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_1_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(SimpleBusCrossbarNto1_1_io_in_2_req_ready),
    .io_in_2_req_valid(SimpleBusCrossbarNto1_1_io_in_2_req_valid),
    .io_in_2_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(SimpleBusCrossbarNto1_1_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(SimpleBusCrossbarNto1_1_io_in_3_req_ready),
    .io_in_3_req_valid(SimpleBusCrossbarNto1_1_io_in_3_req_valid),
    .io_in_3_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr),
    .io_in_3_req_bits_size(SimpleBusCrossbarNto1_1_io_in_3_req_bits_size),
    .io_in_3_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd),
    .io_in_3_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata),
    .io_in_3_resp_ready(SimpleBusCrossbarNto1_1_io_in_3_resp_ready),
    .io_in_3_resp_valid(SimpleBusCrossbarNto1_1_io_in_3_resp_valid),
    .io_in_3_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd),
    .io_in_3_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata)
  );
  EmbeddedTLB EmbeddedTLB ( // @[EmbeddedTLB.scala 421:23]
    .clock(EmbeddedTLB_clock),
    .reset(EmbeddedTLB_reset),
    .io_in_req_ready(EmbeddedTLB_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_io_in_req_bits_addr),
    .io_in_req_bits_user(EmbeddedTLB_io_in_req_bits_user),
    .io_in_resp_ready(EmbeddedTLB_io_in_resp_ready),
    .io_in_resp_valid(EmbeddedTLB_io_in_resp_valid),
    .io_in_resp_bits_rdata(EmbeddedTLB_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(EmbeddedTLB_io_in_resp_bits_user),
    .io_out_req_ready(EmbeddedTLB_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_io_out_req_bits_addr),
    .io_out_req_bits_user(EmbeddedTLB_io_out_req_bits_user),
    .io_out_resp_ready(EmbeddedTLB_io_out_resp_ready),
    .io_out_resp_valid(EmbeddedTLB_io_out_resp_valid),
    .io_out_resp_bits_rdata(EmbeddedTLB_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(EmbeddedTLB_io_out_resp_bits_user),
    .io_mem_req_ready(EmbeddedTLB_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(EmbeddedTLB_io_mem_resp_bits_rdata),
    .io_flush(EmbeddedTLB_io_flush),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_io_csrMMU_priviledgeMode),
    .io_cacheEmpty(EmbeddedTLB_io_cacheEmpty),
    .io_ipf(EmbeddedTLB_io_ipf),
    .CSRSATP(EmbeddedTLB_CSRSATP),
    .MOUFlushTLB(EmbeddedTLB_MOUFlushTLB)
  );
  Cache Cache ( // @[Cache.scala 670:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_user(Cache_io_in_req_bits_user),
    .io_in_resp_ready(Cache_io_in_resp_ready),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(Cache_io_in_resp_bits_user),
    .io_flush(Cache_io_flush),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(Cache_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_io_mmio_req_bits_addr),
    .io_mmio_resp_valid(Cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_io_mmio_resp_bits_rdata),
    .io_empty(Cache_io_empty),
    .MOUFlushICache(Cache_MOUFlushICache)
  );
  EmbeddedTLB_1 EmbeddedTLB_1 ( // @[EmbeddedTLB.scala 421:23]
    .clock(EmbeddedTLB_1_clock),
    .reset(EmbeddedTLB_1_reset),
    .io_in_req_ready(EmbeddedTLB_1_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_1_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_1_io_in_req_bits_addr),
    .io_in_req_bits_size(EmbeddedTLB_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(EmbeddedTLB_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(EmbeddedTLB_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(EmbeddedTLB_1_io_in_req_bits_wdata),
    .io_in_resp_valid(EmbeddedTLB_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(EmbeddedTLB_1_io_in_resp_bits_rdata),
    .io_out_req_ready(EmbeddedTLB_1_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_1_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_1_io_out_req_bits_addr),
    .io_out_req_bits_size(EmbeddedTLB_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(EmbeddedTLB_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(EmbeddedTLB_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(EmbeddedTLB_1_io_out_req_bits_wdata),
    .io_out_resp_valid(EmbeddedTLB_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(EmbeddedTLB_1_io_out_resp_bits_rdata),
    .io_mem_req_ready(EmbeddedTLB_1_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_1_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_1_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_1_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_1_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_1_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(EmbeddedTLB_1_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_1_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(EmbeddedTLB_1_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(EmbeddedTLB_1_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(EmbeddedTLB_1_io_csrMMU_loadPF),
    .io_csrMMU_storePF(EmbeddedTLB_1_io_csrMMU_storePF),
    .io_csrMMU_addr(EmbeddedTLB_1_io_csrMMU_addr),
    ._T_28_0(EmbeddedTLB_1__T_28_0),
    .CSRSATP(EmbeddedTLB_1_CSRSATP),
    .amoReq(EmbeddedTLB_1_amoReq),
    .vmEnable_0(EmbeddedTLB_1_vmEnable_0),
    ._T_27_0(EmbeddedTLB_1__T_27_0),
    .MOUFlushTLB(EmbeddedTLB_1_MOUFlushTLB)
  );
  Cache_1 Cache_1 ( // @[Cache.scala 670:35]
    .clock(Cache_1_clock),
    .reset(Cache_1_reset),
    .io_in_req_ready(Cache_1_io_in_req_ready),
    .io_in_req_valid(Cache_1_io_in_req_valid),
    .io_in_req_bits_addr(Cache_1_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_1_io_in_req_bits_wdata),
    .io_in_resp_ready(Cache_1_io_in_resp_ready),
    .io_in_resp_valid(Cache_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_1_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_1_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_1_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_1_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_1_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_1_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_1_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_1_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_1_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(Cache_1_io_out_coh_req_ready),
    .io_out_coh_req_valid(Cache_1_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(Cache_1_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(Cache_1_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_valid(Cache_1_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(Cache_1_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(Cache_1_io_out_coh_resp_bits_rdata),
    .io_mmio_req_ready(Cache_1_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_1_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_1_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(Cache_1_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(Cache_1_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(Cache_1_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(Cache_1_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(Cache_1_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_1_io_mmio_resp_bits_rdata)
  );
  assign io_imem_mem_req_valid = Cache_io_out_mem_req_valid; // @[NutCore.scala 156:13]
  assign io_imem_mem_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutCore.scala 156:13]
  assign io_imem_mem_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutCore.scala 156:13]
  assign io_imem_mem_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutCore.scala 156:13]
  assign io_dmem_mem_req_valid = Cache_1_io_out_mem_req_valid; // @[NutCore.scala 161:13]
  assign io_dmem_mem_req_bits_addr = Cache_1_io_out_mem_req_bits_addr; // @[NutCore.scala 161:13]
  assign io_dmem_mem_req_bits_cmd = Cache_1_io_out_mem_req_bits_cmd; // @[NutCore.scala 161:13]
  assign io_dmem_mem_req_bits_wdata = Cache_1_io_out_mem_req_bits_wdata; // @[NutCore.scala 161:13]
  assign io_dmem_coh_req_ready = Cache_1_io_out_coh_req_ready; // @[NutCore.scala 161:13]
  assign io_dmem_coh_resp_valid = Cache_1_io_out_coh_resp_valid; // @[NutCore.scala 161:13]
  assign io_dmem_coh_resp_bits_cmd = Cache_1_io_out_coh_resp_bits_cmd; // @[NutCore.scala 161:13]
  assign io_dmem_coh_resp_bits_rdata = Cache_1_io_out_coh_resp_bits_rdata; // @[NutCore.scala 161:13]
  assign io_mmio_req_valid = SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 170:13]
  assign io_mmio_req_bits_addr = SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 170:13]
  assign io_mmio_req_bits_size = SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 170:13]
  assign io_mmio_req_bits_cmd = SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 170:13]
  assign io_mmio_req_bits_wmask = SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 170:13]
  assign io_mmio_req_bits_wdata = SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 170:13]
  assign io_frontend_req_ready = SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 168:23]
  assign io_frontend_resp_valid = SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 168:23]
  assign io_frontend_resp_bits_cmd = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 168:23]
  assign io_frontend_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 168:23]
  assign perfCnts_2 = Backend_inorder_perfCnts_2;
  assign io_in_bits_decode_cf_pc = Backend_inorder_io_in_bits_decode_cf_pc;
  assign io_wb_rfDest = Backend_inorder_io_wb_rfDest;
  assign io_wb_rfWen = Backend_inorder_io_wb_rfWen;
  assign io_wb_rfData = Backend_inorder_io_wb_rfData;
  assign io_in_valid_0 = Backend_inorder_io_in_valid_0;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_imem_req_ready = EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 422:17]
  assign frontend_io_imem_resp_valid = EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 422:17]
  assign frontend_io_imem_resp_bits_rdata = EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 422:17]
  assign frontend_io_imem_resp_bits_user = EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 422:17]
  assign frontend_io_out_0_ready = _T_9 | ~frontend_io_out_0_valid; // @[PipelineVector.scala 50:36]
  assign frontend_io_out_1_ready = _T_9 | ~frontend_io_out_1_valid; // @[PipelineVector.scala 51:36]
  assign frontend_io_redirect_target = Backend_inorder_io_redirect_target; // @[NutCore.scala 164:26]
  assign frontend_io_redirect_valid = Backend_inorder_io_redirect_valid; // @[NutCore.scala 164:26]
  assign frontend_io_ipf = EmbeddedTLB_io_ipf; // @[NutCore.scala 155:21]
  assign frontend_flushICache = Backend_inorder_flushICache;
  assign frontend_REG_0_valid = Backend_inorder_REG_0_valid;
  assign frontend_REG_0_pc = Backend_inorder_REG_0_pc;
  assign frontend_REG_0_isMissPredict = Backend_inorder_REG_0_isMissPredict;
  assign frontend_REG_0_actualTarget = Backend_inorder_REG_0_actualTarget;
  assign frontend_REG_0_actualTaken = Backend_inorder_REG_0_actualTaken;
  assign frontend_REG_0_fuOpType = Backend_inorder_REG_0_fuOpType;
  assign frontend_REG_0_btbType = Backend_inorder_REG_0_btbType;
  assign frontend_REG_0_isRVC = Backend_inorder_REG_0_isRVC;
  assign frontend_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign frontend_intrVec = Backend_inorder_intrVec;
  assign frontend_flushTLB = Backend_inorder_flushTLB;
  assign Backend_inorder_clock = clock;
  assign Backend_inorder_reset = reset;
  assign Backend_inorder_io_in_0_valid = REG_1 != REG_2; // @[PipelineVector.scala 56:34]
  assign Backend_inorder_io_in_0_bits_cf_instr = 2'h3 == REG_2 ? REG__3_cf_instr : _GEN_1415; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_pc = 2'h3 == REG_2 ? REG__3_cf_pc : _GEN_1411; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_pnpc = 2'h3 == REG_2 ? REG__3_cf_pnpc : _GEN_1407; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == REG_2 ? REG__3_cf_exceptionVec_1 : _GEN_1335; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == REG_2 ? REG__3_cf_exceptionVec_2 : _GEN_1339; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == REG_2 ? REG__3_cf_exceptionVec_12 : _GEN_1379; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_0 = 2'h3 == REG_2 ? REG__3_cf_intrVec_0 : _GEN_1283; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_1 = 2'h3 == REG_2 ? REG__3_cf_intrVec_1 : _GEN_1287; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_2 = 2'h3 == REG_2 ? REG__3_cf_intrVec_2 : _GEN_1291; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_3 = 2'h3 == REG_2 ? REG__3_cf_intrVec_3 : _GEN_1295; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_4 = 2'h3 == REG_2 ? REG__3_cf_intrVec_4 : _GEN_1299; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_5 = 2'h3 == REG_2 ? REG__3_cf_intrVec_5 : _GEN_1303; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_6 = 2'h3 == REG_2 ? REG__3_cf_intrVec_6 : _GEN_1307; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_7 = 2'h3 == REG_2 ? REG__3_cf_intrVec_7 : _GEN_1311; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_8 = 2'h3 == REG_2 ? REG__3_cf_intrVec_8 : _GEN_1315; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_9 = 2'h3 == REG_2 ? REG__3_cf_intrVec_9 : _GEN_1319; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_10 = 2'h3 == REG_2 ? REG__3_cf_intrVec_10 : _GEN_1323; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_11 = 2'h3 == REG_2 ? REG__3_cf_intrVec_11 : _GEN_1327; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_brIdx = 2'h3 == REG_2 ? REG__3_cf_brIdx : _GEN_1279; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_crossPageIPFFix = 2'h3 == REG_2 ? REG__3_cf_crossPageIPFFix : _GEN_1271; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_cf_runahead_checkpoint_id = 2'h3 == REG_2 ? REG__3_cf_runahead_checkpoint_id :
    _GEN_1267; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_src1Type = 2'h3 == REG_2 ? REG__3_ctrl_src1Type : _GEN_1259; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_src2Type = 2'h3 == REG_2 ? REG__3_ctrl_src2Type : _GEN_1255; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_fuType = 2'h3 == REG_2 ? REG__3_ctrl_fuType : _GEN_1251; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_fuOpType = 2'h3 == REG_2 ? REG__3_ctrl_fuOpType : _GEN_1247; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == REG_2 ? REG__3_ctrl_rfSrc1 : _GEN_1243; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == REG_2 ? REG__3_ctrl_rfSrc2 : _GEN_1239; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_rfWen = 2'h3 == REG_2 ? REG__3_ctrl_rfWen : _GEN_1235; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_rfDest = 2'h3 == REG_2 ? REG__3_ctrl_rfDest : _GEN_1231; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_vtag = 2'h3 == REG_2 ? REG__3_ctrl_vtag : _GEN_1207; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_vec_addr = 2'h3 == REG_2 ? REG__3_ctrl_vec_addr : _GEN_1203; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_length_k = 2'h3 == REG_2 ? REG__3_ctrl_length_k : _GEN_1199; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_ctrl_algorithm = 2'h3 == REG_2 ? REG__3_ctrl_algorithm : _GEN_1195; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_in_0_bits_data_imm = 2'h3 == REG_2 ? REG__3_data_imm : _GEN_1183; // @[PipelineVector.scala 55:{15,15}]
  assign Backend_inorder_io_flush = frontend_io_flushVec[3:2]; // @[NutCore.scala 165:45]
  assign Backend_inorder_io_dmem_req_ready = EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 422:17]
  assign Backend_inorder_io_dmem_resp_valid = EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 422:17]
  assign Backend_inorder_io_dmem_resp_bits_rdata = EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 422:17]
  assign Backend_inorder_io_memMMU_dmem_loadPF = EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 425:21]
  assign Backend_inorder_io_memMMU_dmem_storePF = EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 425:21]
  assign Backend_inorder_io_memMMU_dmem_addr = EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 425:21]
  assign Backend_inorder__T_28 = EmbeddedTLB_1__T_28_0;
  assign Backend_inorder_io_extra_mtip = io_extra_mtip;
  assign Backend_inorder_io_extra_meip_0 = io_extra_meip_0;
  assign Backend_inorder_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign Backend_inorder__T_27 = EmbeddedTLB_1__T_27_0;
  assign Backend_inorder_io_extra_msip = io_extra_msip;
  assign SimpleBusCrossbarNto1_clock = clock;
  assign SimpleBusCrossbarNto1_reset = reset;
  assign SimpleBusCrossbarNto1_io_in_0_req_valid = Cache_io_mmio_req_valid; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_addr = Cache_io_mmio_req_bits_addr; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_cmd = 4'h0; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wmask = 8'h0; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wdata = 64'h0; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_valid = Cache_1_io_mmio_req_valid; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_addr = Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_size = Cache_1_io_mmio_req_bits_size; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_cmd = Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wmask = Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wdata = Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 677:13]
  assign SimpleBusCrossbarNto1_io_out_req_ready = io_mmio_req_ready; // @[NutCore.scala 170:13]
  assign SimpleBusCrossbarNto1_io_out_resp_valid = io_mmio_resp_valid; // @[NutCore.scala 170:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[NutCore.scala 170:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[NutCore.scala 170:13]
  assign SimpleBusCrossbarNto1_1_clock = clock;
  assign SimpleBusCrossbarNto1_1_reset = reset;
  assign SimpleBusCrossbarNto1_1_io_in_0_req_valid = EmbeddedTLB_1_io_out_req_valid; // @[NutCore.scala 160:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr = EmbeddedTLB_1_io_out_req_bits_addr; // @[NutCore.scala 160:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_size = EmbeddedTLB_1_io_out_req_bits_size; // @[NutCore.scala 160:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd = EmbeddedTLB_1_io_out_req_bits_cmd; // @[NutCore.scala 160:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask = EmbeddedTLB_1_io_out_req_bits_wmask; // @[NutCore.scala 160:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata = EmbeddedTLB_1_io_out_req_bits_wdata; // @[NutCore.scala 160:23]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_valid = EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr = EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd = EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata = EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_valid = EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr = EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd = EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata = EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 423:18]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_valid = io_frontend_req_valid; // @[NutCore.scala 168:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr = io_frontend_req_bits_addr; // @[NutCore.scala 168:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_size = io_frontend_req_bits_size; // @[NutCore.scala 168:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd = io_frontend_req_bits_cmd; // @[NutCore.scala 168:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask = io_frontend_req_bits_wmask; // @[NutCore.scala 168:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata = io_frontend_req_bits_wdata; // @[NutCore.scala 168:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_resp_ready = io_frontend_resp_ready; // @[NutCore.scala 168:23]
  assign SimpleBusCrossbarNto1_1_io_out_req_ready = Cache_1_io_in_req_ready; // @[Cache.scala 676:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_valid = Cache_1_io_in_resp_valid; // @[Cache.scala 676:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd = Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 676:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata = Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 676:17]
  assign EmbeddedTLB_clock = clock;
  assign EmbeddedTLB_reset = reset;
  assign EmbeddedTLB_io_in_req_valid = frontend_io_imem_req_valid; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_io_in_resp_ready = frontend_io_imem_resp_ready; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_io_out_req_ready = Cache_io_in_req_ready; // @[Cache.scala 676:17]
  assign EmbeddedTLB_io_out_resp_valid = Cache_io_in_resp_valid; // @[Cache.scala 676:17]
  assign EmbeddedTLB_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[Cache.scala 676:17]
  assign EmbeddedTLB_io_out_resp_bits_user = Cache_io_in_resp_bits_user; // @[Cache.scala 676:17]
  assign EmbeddedTLB_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[EmbeddedTLB.scala 423:18]
  assign EmbeddedTLB_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[EmbeddedTLB.scala 423:18]
  assign EmbeddedTLB_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[EmbeddedTLB.scala 423:18]
  assign EmbeddedTLB_io_flush = frontend_io_flushVec[0]; // @[NutCore.scala 154:104]
  assign EmbeddedTLB_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_imem_priviledgeMode; // @[EmbeddedTLB.scala 425:21]
  assign EmbeddedTLB_io_cacheEmpty = Cache_io_empty; // @[Cache.scala 678:11]
  assign EmbeddedTLB_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = EmbeddedTLB_io_out_req_valid; // @[Cache.scala 676:17]
  assign Cache_io_in_req_bits_addr = EmbeddedTLB_io_out_req_bits_addr; // @[Cache.scala 676:17]
  assign Cache_io_in_req_bits_user = EmbeddedTLB_io_out_req_bits_user; // @[Cache.scala 676:17]
  assign Cache_io_in_resp_ready = EmbeddedTLB_io_out_resp_ready; // @[Cache.scala 676:17]
  assign Cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign Cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[NutCore.scala 156:13]
  assign Cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[NutCore.scala 156:13]
  assign Cache_io_out_mem_resp_bits_cmd = io_imem_mem_resp_bits_cmd; // @[NutCore.scala 156:13]
  assign Cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[NutCore.scala 156:13]
  assign Cache_io_mmio_req_ready = SimpleBusCrossbarNto1_io_in_0_req_ready; // @[Cache.scala 677:13]
  assign Cache_io_mmio_resp_valid = SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[Cache.scala 677:13]
  assign Cache_io_mmio_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[Cache.scala 677:13]
  assign Cache_MOUFlushICache = Backend_inorder_flushICache;
  assign EmbeddedTLB_1_clock = clock;
  assign EmbeddedTLB_1_reset = reset;
  assign EmbeddedTLB_1_io_in_req_valid = Backend_inorder_io_dmem_req_valid; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_1_io_in_req_bits_addr = Backend_inorder_io_dmem_req_bits_addr; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_1_io_in_req_bits_size = Backend_inorder_io_dmem_req_bits_size; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_1_io_in_req_bits_cmd = Backend_inorder_io_dmem_req_bits_cmd; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_1_io_in_req_bits_wmask = Backend_inorder_io_dmem_req_bits_wmask; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_1_io_in_req_bits_wdata = Backend_inorder_io_dmem_req_bits_wdata; // @[EmbeddedTLB.scala 422:17]
  assign EmbeddedTLB_1_io_out_req_ready = SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 160:23]
  assign EmbeddedTLB_1_io_out_resp_valid = SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 160:23]
  assign EmbeddedTLB_1_io_out_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 160:23]
  assign EmbeddedTLB_1_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[EmbeddedTLB.scala 423:18]
  assign EmbeddedTLB_1_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[EmbeddedTLB.scala 423:18]
  assign EmbeddedTLB_1_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[EmbeddedTLB.scala 423:18]
  assign EmbeddedTLB_1_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[EmbeddedTLB.scala 425:21]
  assign EmbeddedTLB_1_io_csrMMU_status_sum = Backend_inorder_io_memMMU_dmem_status_sum; // @[EmbeddedTLB.scala 425:21]
  assign EmbeddedTLB_1_io_csrMMU_status_mxr = Backend_inorder_io_memMMU_dmem_status_mxr; // @[EmbeddedTLB.scala 425:21]
  assign EmbeddedTLB_1_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_1_amoReq = Backend_inorder_amoReq;
  assign EmbeddedTLB_1_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_1_clock = clock;
  assign Cache_1_reset = reset;
  assign Cache_1_io_in_req_valid = SimpleBusCrossbarNto1_1_io_out_req_valid; // @[Cache.scala 676:17]
  assign Cache_1_io_in_req_bits_addr = SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[Cache.scala 676:17]
  assign Cache_1_io_in_req_bits_size = SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[Cache.scala 676:17]
  assign Cache_1_io_in_req_bits_cmd = SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[Cache.scala 676:17]
  assign Cache_1_io_in_req_bits_wmask = SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[Cache.scala 676:17]
  assign Cache_1_io_in_req_bits_wdata = SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[Cache.scala 676:17]
  assign Cache_1_io_in_resp_ready = SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[Cache.scala 676:17]
  assign Cache_1_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[NutCore.scala 161:13]
  assign Cache_1_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[NutCore.scala 161:13]
  assign Cache_1_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[NutCore.scala 161:13]
  assign Cache_1_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[NutCore.scala 161:13]
  assign Cache_1_io_out_coh_req_valid = io_dmem_coh_req_valid; // @[NutCore.scala 161:13]
  assign Cache_1_io_out_coh_req_bits_addr = io_dmem_coh_req_bits_addr; // @[NutCore.scala 161:13]
  assign Cache_1_io_out_coh_req_bits_wdata = io_dmem_coh_req_bits_wdata; // @[NutCore.scala 161:13]
  assign Cache_1_io_mmio_req_ready = SimpleBusCrossbarNto1_io_in_1_req_ready; // @[Cache.scala 677:13]
  assign Cache_1_io_mmio_resp_valid = SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[Cache.scala 677:13]
  assign Cache_1_io_mmio_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[Cache.scala 677:13]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_instr <= _GEN_468;
        end
      end else begin
        REG__0_cf_instr <= _GEN_468;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_pc <= _GEN_464;
        end
      end else begin
        REG__0_cf_pc <= _GEN_464;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_pnpc <= _GEN_460;
        end
      end else begin
        REG__0_cf_pnpc <= _GEN_460;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_1 <= _GEN_388;
        end
      end else begin
        REG__0_cf_exceptionVec_1 <= _GEN_388;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_2 <= _GEN_392;
        end
      end else begin
        REG__0_cf_exceptionVec_2 <= _GEN_392;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_12 <= _GEN_432;
        end
      end else begin
        REG__0_cf_exceptionVec_12 <= _GEN_432;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_0 <= _GEN_336;
        end
      end else begin
        REG__0_cf_intrVec_0 <= _GEN_336;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_1 <= _GEN_340;
        end
      end else begin
        REG__0_cf_intrVec_1 <= _GEN_340;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_2 <= _GEN_344;
        end
      end else begin
        REG__0_cf_intrVec_2 <= _GEN_344;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_3 <= _GEN_348;
        end
      end else begin
        REG__0_cf_intrVec_3 <= _GEN_348;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_4 <= _GEN_352;
        end
      end else begin
        REG__0_cf_intrVec_4 <= _GEN_352;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_5 <= _GEN_356;
        end
      end else begin
        REG__0_cf_intrVec_5 <= _GEN_356;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_6 <= _GEN_360;
        end
      end else begin
        REG__0_cf_intrVec_6 <= _GEN_360;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_7 <= _GEN_364;
        end
      end else begin
        REG__0_cf_intrVec_7 <= _GEN_364;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_8 <= _GEN_368;
        end
      end else begin
        REG__0_cf_intrVec_8 <= _GEN_368;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_9 <= _GEN_372;
        end
      end else begin
        REG__0_cf_intrVec_9 <= _GEN_372;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_10 <= _GEN_376;
        end
      end else begin
        REG__0_cf_intrVec_10 <= _GEN_376;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_11 <= _GEN_380;
        end
      end else begin
        REG__0_cf_intrVec_11 <= _GEN_380;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_brIdx <= _GEN_332;
        end
      end else begin
        REG__0_cf_brIdx <= _GEN_332;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_crossPageIPFFix <= _GEN_324;
        end
      end else begin
        REG__0_cf_crossPageIPFFix <= _GEN_324;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_runahead_checkpoint_id <= _GEN_320;
        end
      end else begin
        REG__0_cf_runahead_checkpoint_id <= _GEN_320;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_src1Type <= _GEN_312;
        end
      end else begin
        REG__0_ctrl_src1Type <= _GEN_312;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_src2Type <= _GEN_308;
        end
      end else begin
        REG__0_ctrl_src2Type <= _GEN_308;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_fuType <= _GEN_304;
        end
      end else begin
        REG__0_ctrl_fuType <= _GEN_304;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_fuOpType <= _GEN_300;
        end
      end else begin
        REG__0_ctrl_fuOpType <= _GEN_300;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfSrc1 <= _GEN_296;
        end
      end else begin
        REG__0_ctrl_rfSrc1 <= _GEN_296;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfSrc2 <= _GEN_292;
        end
      end else begin
        REG__0_ctrl_rfSrc2 <= _GEN_292;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfWen <= _GEN_288;
        end
      end else begin
        REG__0_ctrl_rfWen <= _GEN_288;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfDest <= _GEN_284;
        end
      end else begin
        REG__0_ctrl_rfDest <= _GEN_284;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_vtag <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_vtag <= _REG_T_20_ctrl_vtag; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_vtag <= _GEN_260;
        end
      end else begin
        REG__0_ctrl_vtag <= _GEN_260;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_vec_addr <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_vec_addr <= _REG_T_20_ctrl_vec_addr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_vec_addr <= _GEN_256;
        end
      end else begin
        REG__0_ctrl_vec_addr <= _GEN_256;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_length_k <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_length_k <= _REG_T_20_ctrl_length_k; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_length_k <= _GEN_252;
        end
      end else begin
        REG__0_ctrl_length_k <= _GEN_252;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_algorithm <= 2'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_algorithm <= _REG_T_20_ctrl_algorithm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_algorithm <= _GEN_248;
        end
      end else begin
        REG__0_ctrl_algorithm <= _GEN_248;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_data_imm <= _GEN_236;
        end
      end else begin
        REG__0_data_imm <= _GEN_236;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_instr <= _GEN_469;
        end
      end else begin
        REG__1_cf_instr <= _GEN_469;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_pc <= _GEN_465;
        end
      end else begin
        REG__1_cf_pc <= _GEN_465;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_pnpc <= _GEN_461;
        end
      end else begin
        REG__1_cf_pnpc <= _GEN_461;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_1 <= _GEN_389;
        end
      end else begin
        REG__1_cf_exceptionVec_1 <= _GEN_389;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_2 <= _GEN_393;
        end
      end else begin
        REG__1_cf_exceptionVec_2 <= _GEN_393;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_12 <= _GEN_433;
        end
      end else begin
        REG__1_cf_exceptionVec_12 <= _GEN_433;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_0 <= _GEN_337;
        end
      end else begin
        REG__1_cf_intrVec_0 <= _GEN_337;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_1 <= _GEN_341;
        end
      end else begin
        REG__1_cf_intrVec_1 <= _GEN_341;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_2 <= _GEN_345;
        end
      end else begin
        REG__1_cf_intrVec_2 <= _GEN_345;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_3 <= _GEN_349;
        end
      end else begin
        REG__1_cf_intrVec_3 <= _GEN_349;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_4 <= _GEN_353;
        end
      end else begin
        REG__1_cf_intrVec_4 <= _GEN_353;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_5 <= _GEN_357;
        end
      end else begin
        REG__1_cf_intrVec_5 <= _GEN_357;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_6 <= _GEN_361;
        end
      end else begin
        REG__1_cf_intrVec_6 <= _GEN_361;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_7 <= _GEN_365;
        end
      end else begin
        REG__1_cf_intrVec_7 <= _GEN_365;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_8 <= _GEN_369;
        end
      end else begin
        REG__1_cf_intrVec_8 <= _GEN_369;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_9 <= _GEN_373;
        end
      end else begin
        REG__1_cf_intrVec_9 <= _GEN_373;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_10 <= _GEN_377;
        end
      end else begin
        REG__1_cf_intrVec_10 <= _GEN_377;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_11 <= _GEN_381;
        end
      end else begin
        REG__1_cf_intrVec_11 <= _GEN_381;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_brIdx <= _GEN_333;
        end
      end else begin
        REG__1_cf_brIdx <= _GEN_333;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_crossPageIPFFix <= _GEN_325;
        end
      end else begin
        REG__1_cf_crossPageIPFFix <= _GEN_325;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_runahead_checkpoint_id <= _GEN_321;
        end
      end else begin
        REG__1_cf_runahead_checkpoint_id <= _GEN_321;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_src1Type <= _GEN_313;
        end
      end else begin
        REG__1_ctrl_src1Type <= _GEN_313;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_src2Type <= _GEN_309;
        end
      end else begin
        REG__1_ctrl_src2Type <= _GEN_309;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_fuType <= _GEN_305;
        end
      end else begin
        REG__1_ctrl_fuType <= _GEN_305;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_fuOpType <= _GEN_301;
        end
      end else begin
        REG__1_ctrl_fuOpType <= _GEN_301;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfSrc1 <= _GEN_297;
        end
      end else begin
        REG__1_ctrl_rfSrc1 <= _GEN_297;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfSrc2 <= _GEN_293;
        end
      end else begin
        REG__1_ctrl_rfSrc2 <= _GEN_293;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfWen <= _GEN_289;
        end
      end else begin
        REG__1_ctrl_rfWen <= _GEN_289;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfDest <= _GEN_285;
        end
      end else begin
        REG__1_ctrl_rfDest <= _GEN_285;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_vtag <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_vtag <= _REG_T_20_ctrl_vtag; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_vtag <= _GEN_261;
        end
      end else begin
        REG__1_ctrl_vtag <= _GEN_261;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_vec_addr <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_vec_addr <= _REG_T_20_ctrl_vec_addr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_vec_addr <= _GEN_257;
        end
      end else begin
        REG__1_ctrl_vec_addr <= _GEN_257;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_length_k <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_length_k <= _REG_T_20_ctrl_length_k; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_length_k <= _GEN_253;
        end
      end else begin
        REG__1_ctrl_length_k <= _GEN_253;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_algorithm <= 2'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_algorithm <= _REG_T_20_ctrl_algorithm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_algorithm <= _GEN_249;
        end
      end else begin
        REG__1_ctrl_algorithm <= _GEN_249;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_data_imm <= _GEN_237;
        end
      end else begin
        REG__1_data_imm <= _GEN_237;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_instr <= _GEN_470;
        end
      end else begin
        REG__2_cf_instr <= _GEN_470;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_pc <= _GEN_466;
        end
      end else begin
        REG__2_cf_pc <= _GEN_466;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_pnpc <= _GEN_462;
        end
      end else begin
        REG__2_cf_pnpc <= _GEN_462;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_1 <= _GEN_390;
        end
      end else begin
        REG__2_cf_exceptionVec_1 <= _GEN_390;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_2 <= _GEN_394;
        end
      end else begin
        REG__2_cf_exceptionVec_2 <= _GEN_394;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_12 <= _GEN_434;
        end
      end else begin
        REG__2_cf_exceptionVec_12 <= _GEN_434;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_0 <= _GEN_338;
        end
      end else begin
        REG__2_cf_intrVec_0 <= _GEN_338;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_1 <= _GEN_342;
        end
      end else begin
        REG__2_cf_intrVec_1 <= _GEN_342;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_2 <= _GEN_346;
        end
      end else begin
        REG__2_cf_intrVec_2 <= _GEN_346;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_3 <= _GEN_350;
        end
      end else begin
        REG__2_cf_intrVec_3 <= _GEN_350;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_4 <= _GEN_354;
        end
      end else begin
        REG__2_cf_intrVec_4 <= _GEN_354;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_5 <= _GEN_358;
        end
      end else begin
        REG__2_cf_intrVec_5 <= _GEN_358;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_6 <= _GEN_362;
        end
      end else begin
        REG__2_cf_intrVec_6 <= _GEN_362;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_7 <= _GEN_366;
        end
      end else begin
        REG__2_cf_intrVec_7 <= _GEN_366;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_8 <= _GEN_370;
        end
      end else begin
        REG__2_cf_intrVec_8 <= _GEN_370;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_9 <= _GEN_374;
        end
      end else begin
        REG__2_cf_intrVec_9 <= _GEN_374;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_10 <= _GEN_378;
        end
      end else begin
        REG__2_cf_intrVec_10 <= _GEN_378;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_11 <= _GEN_382;
        end
      end else begin
        REG__2_cf_intrVec_11 <= _GEN_382;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_brIdx <= _GEN_334;
        end
      end else begin
        REG__2_cf_brIdx <= _GEN_334;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_crossPageIPFFix <= _GEN_326;
        end
      end else begin
        REG__2_cf_crossPageIPFFix <= _GEN_326;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_runahead_checkpoint_id <= _GEN_322;
        end
      end else begin
        REG__2_cf_runahead_checkpoint_id <= _GEN_322;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_src1Type <= _GEN_314;
        end
      end else begin
        REG__2_ctrl_src1Type <= _GEN_314;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_src2Type <= _GEN_310;
        end
      end else begin
        REG__2_ctrl_src2Type <= _GEN_310;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_fuType <= _GEN_306;
        end
      end else begin
        REG__2_ctrl_fuType <= _GEN_306;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_fuOpType <= _GEN_302;
        end
      end else begin
        REG__2_ctrl_fuOpType <= _GEN_302;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfSrc1 <= _GEN_298;
        end
      end else begin
        REG__2_ctrl_rfSrc1 <= _GEN_298;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfSrc2 <= _GEN_294;
        end
      end else begin
        REG__2_ctrl_rfSrc2 <= _GEN_294;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfWen <= _GEN_290;
        end
      end else begin
        REG__2_ctrl_rfWen <= _GEN_290;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfDest <= _GEN_286;
        end
      end else begin
        REG__2_ctrl_rfDest <= _GEN_286;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_vtag <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_vtag <= _REG_T_20_ctrl_vtag; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_vtag <= _GEN_262;
        end
      end else begin
        REG__2_ctrl_vtag <= _GEN_262;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_vec_addr <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_vec_addr <= _REG_T_20_ctrl_vec_addr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_vec_addr <= _GEN_258;
        end
      end else begin
        REG__2_ctrl_vec_addr <= _GEN_258;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_length_k <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_length_k <= _REG_T_20_ctrl_length_k; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_length_k <= _GEN_254;
        end
      end else begin
        REG__2_ctrl_length_k <= _GEN_254;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_algorithm <= 2'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_algorithm <= _REG_T_20_ctrl_algorithm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_algorithm <= _GEN_250;
        end
      end else begin
        REG__2_ctrl_algorithm <= _GEN_250;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_data_imm <= _GEN_238;
        end
      end else begin
        REG__2_data_imm <= _GEN_238;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_instr <= _GEN_471;
        end
      end else begin
        REG__3_cf_instr <= _GEN_471;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_pc <= _GEN_467;
        end
      end else begin
        REG__3_cf_pc <= _GEN_467;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_pnpc <= _GEN_463;
        end
      end else begin
        REG__3_cf_pnpc <= _GEN_463;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_1 <= _GEN_391;
        end
      end else begin
        REG__3_cf_exceptionVec_1 <= _GEN_391;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_2 <= _GEN_395;
        end
      end else begin
        REG__3_cf_exceptionVec_2 <= _GEN_395;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_12 <= _GEN_435;
        end
      end else begin
        REG__3_cf_exceptionVec_12 <= _GEN_435;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_0 <= _GEN_339;
        end
      end else begin
        REG__3_cf_intrVec_0 <= _GEN_339;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_1 <= _GEN_343;
        end
      end else begin
        REG__3_cf_intrVec_1 <= _GEN_343;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_2 <= _GEN_347;
        end
      end else begin
        REG__3_cf_intrVec_2 <= _GEN_347;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_3 <= _GEN_351;
        end
      end else begin
        REG__3_cf_intrVec_3 <= _GEN_351;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_4 <= _GEN_355;
        end
      end else begin
        REG__3_cf_intrVec_4 <= _GEN_355;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_5 <= _GEN_359;
        end
      end else begin
        REG__3_cf_intrVec_5 <= _GEN_359;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_6 <= _GEN_363;
        end
      end else begin
        REG__3_cf_intrVec_6 <= _GEN_363;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_7 <= _GEN_367;
        end
      end else begin
        REG__3_cf_intrVec_7 <= _GEN_367;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_8 <= _GEN_371;
        end
      end else begin
        REG__3_cf_intrVec_8 <= _GEN_371;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_9 <= _GEN_375;
        end
      end else begin
        REG__3_cf_intrVec_9 <= _GEN_375;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_10 <= _GEN_379;
        end
      end else begin
        REG__3_cf_intrVec_10 <= _GEN_379;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_11 <= _GEN_383;
        end
      end else begin
        REG__3_cf_intrVec_11 <= _GEN_383;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_brIdx <= _GEN_335;
        end
      end else begin
        REG__3_cf_brIdx <= _GEN_335;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_crossPageIPFFix <= _GEN_327;
        end
      end else begin
        REG__3_cf_crossPageIPFFix <= _GEN_327;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_runahead_checkpoint_id <= 64'h0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_runahead_checkpoint_id <= _GEN_323;
        end
      end else begin
        REG__3_cf_runahead_checkpoint_id <= _GEN_323;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_src1Type <= _GEN_315;
        end
      end else begin
        REG__3_ctrl_src1Type <= _GEN_315;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_src2Type <= _GEN_311;
        end
      end else begin
        REG__3_ctrl_src2Type <= _GEN_311;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_fuType <= _GEN_307;
        end
      end else begin
        REG__3_ctrl_fuType <= _GEN_307;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_fuOpType <= _GEN_303;
        end
      end else begin
        REG__3_ctrl_fuOpType <= _GEN_303;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfSrc1 <= _GEN_299;
        end
      end else begin
        REG__3_ctrl_rfSrc1 <= _GEN_299;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfSrc2 <= _GEN_295;
        end
      end else begin
        REG__3_ctrl_rfSrc2 <= _GEN_295;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfWen <= _GEN_291;
        end
      end else begin
        REG__3_ctrl_rfWen <= _GEN_291;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfDest <= _GEN_287;
        end
      end else begin
        REG__3_ctrl_rfDest <= _GEN_287;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_vtag <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_vtag <= _REG_T_20_ctrl_vtag; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_vtag <= _GEN_263;
        end
      end else begin
        REG__3_ctrl_vtag <= _GEN_263;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_vec_addr <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_vec_addr <= _REG_T_20_ctrl_vec_addr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_vec_addr <= _GEN_259;
        end
      end else begin
        REG__3_ctrl_vec_addr <= _GEN_259;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_length_k <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_length_k <= _REG_T_20_ctrl_length_k; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_length_k <= _GEN_255;
        end
      end else begin
        REG__3_ctrl_length_k <= _GEN_255;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_algorithm <= 2'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_algorithm <= _REG_T_20_ctrl_algorithm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_algorithm <= _GEN_251;
        end
      end else begin
        REG__3_ctrl_algorithm <= _GEN_251;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_data_imm <= _GEN_239;
        end
      end else begin
        REG__3_data_imm <= _GEN_239;
      end
    end
    if (reset) begin // @[PipelineVector.scala 30:33]
      REG_1 <= 2'h0; // @[PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[PipelineVector.scala 71:16]
      REG_1 <= 2'h0; // @[PipelineVector.scala 72:24]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      REG_1 <= _T_22; // @[PipelineVector.scala 47:24]
    end
    if (reset) begin // @[PipelineVector.scala 31:33]
      REG_2 <= 2'h0; // @[PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[PipelineVector.scala 71:16]
      REG_2 <= 2'h0; // @[PipelineVector.scala 73:24]
    end else if (_T_35) begin // @[PipelineVector.scala 66:22]
      REG_2 <= _T_37; // @[PipelineVector.scala 67:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG__0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  REG__0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  REG__0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG__0_cf_intrVec_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG__0_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG__0_cf_intrVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG__0_cf_intrVec_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG__0_cf_intrVec_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG__0_cf_intrVec_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG__0_cf_intrVec_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG__0_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG__0_cf_intrVec_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  REG__0_cf_intrVec_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG__0_cf_intrVec_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG__0_cf_intrVec_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG__0_cf_brIdx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  REG__0_cf_crossPageIPFFix = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  REG__0_cf_runahead_checkpoint_id = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  REG__0_ctrl_src1Type = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  REG__0_ctrl_src2Type = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  REG__0_ctrl_fuType = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  REG__0_ctrl_fuOpType = _RAND_24[6:0];
  _RAND_25 = {1{`RANDOM}};
  REG__0_ctrl_rfSrc1 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  REG__0_ctrl_rfSrc2 = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  REG__0_ctrl_rfWen = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  REG__0_ctrl_rfDest = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  REG__0_ctrl_vtag = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  REG__0_ctrl_vec_addr = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  REG__0_ctrl_length_k = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  REG__0_ctrl_algorithm = _RAND_32[1:0];
  _RAND_33 = {2{`RANDOM}};
  REG__0_data_imm = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  REG__1_cf_instr = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  REG__1_cf_pc = _RAND_35[38:0];
  _RAND_36 = {2{`RANDOM}};
  REG__1_cf_pnpc = _RAND_36[38:0];
  _RAND_37 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_12 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  REG__1_cf_intrVec_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  REG__1_cf_intrVec_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  REG__1_cf_intrVec_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  REG__1_cf_intrVec_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  REG__1_cf_intrVec_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG__1_cf_intrVec_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG__1_cf_intrVec_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  REG__1_cf_intrVec_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG__1_cf_intrVec_8 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG__1_cf_intrVec_9 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG__1_cf_intrVec_10 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG__1_cf_intrVec_11 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  REG__1_cf_brIdx = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  REG__1_cf_crossPageIPFFix = _RAND_53[0:0];
  _RAND_54 = {2{`RANDOM}};
  REG__1_cf_runahead_checkpoint_id = _RAND_54[63:0];
  _RAND_55 = {1{`RANDOM}};
  REG__1_ctrl_src1Type = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  REG__1_ctrl_src2Type = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  REG__1_ctrl_fuType = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  REG__1_ctrl_fuOpType = _RAND_58[6:0];
  _RAND_59 = {1{`RANDOM}};
  REG__1_ctrl_rfSrc1 = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  REG__1_ctrl_rfSrc2 = _RAND_60[4:0];
  _RAND_61 = {1{`RANDOM}};
  REG__1_ctrl_rfWen = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  REG__1_ctrl_rfDest = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  REG__1_ctrl_vtag = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  REG__1_ctrl_vec_addr = _RAND_64[4:0];
  _RAND_65 = {1{`RANDOM}};
  REG__1_ctrl_length_k = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  REG__1_ctrl_algorithm = _RAND_66[1:0];
  _RAND_67 = {2{`RANDOM}};
  REG__1_data_imm = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  REG__2_cf_instr = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  REG__2_cf_pc = _RAND_69[38:0];
  _RAND_70 = {2{`RANDOM}};
  REG__2_cf_pnpc = _RAND_70[38:0];
  _RAND_71 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_1 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_2 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_12 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  REG__2_cf_intrVec_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  REG__2_cf_intrVec_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  REG__2_cf_intrVec_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  REG__2_cf_intrVec_3 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  REG__2_cf_intrVec_4 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  REG__2_cf_intrVec_5 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  REG__2_cf_intrVec_6 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  REG__2_cf_intrVec_7 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  REG__2_cf_intrVec_8 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  REG__2_cf_intrVec_9 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  REG__2_cf_intrVec_10 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  REG__2_cf_intrVec_11 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  REG__2_cf_brIdx = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  REG__2_cf_crossPageIPFFix = _RAND_87[0:0];
  _RAND_88 = {2{`RANDOM}};
  REG__2_cf_runahead_checkpoint_id = _RAND_88[63:0];
  _RAND_89 = {1{`RANDOM}};
  REG__2_ctrl_src1Type = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  REG__2_ctrl_src2Type = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  REG__2_ctrl_fuType = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  REG__2_ctrl_fuOpType = _RAND_92[6:0];
  _RAND_93 = {1{`RANDOM}};
  REG__2_ctrl_rfSrc1 = _RAND_93[4:0];
  _RAND_94 = {1{`RANDOM}};
  REG__2_ctrl_rfSrc2 = _RAND_94[4:0];
  _RAND_95 = {1{`RANDOM}};
  REG__2_ctrl_rfWen = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  REG__2_ctrl_rfDest = _RAND_96[4:0];
  _RAND_97 = {1{`RANDOM}};
  REG__2_ctrl_vtag = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  REG__2_ctrl_vec_addr = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  REG__2_ctrl_length_k = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  REG__2_ctrl_algorithm = _RAND_100[1:0];
  _RAND_101 = {2{`RANDOM}};
  REG__2_data_imm = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  REG__3_cf_instr = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  REG__3_cf_pc = _RAND_103[38:0];
  _RAND_104 = {2{`RANDOM}};
  REG__3_cf_pnpc = _RAND_104[38:0];
  _RAND_105 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_2 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_12 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG__3_cf_intrVec_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG__3_cf_intrVec_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  REG__3_cf_intrVec_2 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  REG__3_cf_intrVec_3 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  REG__3_cf_intrVec_4 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  REG__3_cf_intrVec_5 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  REG__3_cf_intrVec_6 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  REG__3_cf_intrVec_7 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  REG__3_cf_intrVec_8 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG__3_cf_intrVec_9 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  REG__3_cf_intrVec_10 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  REG__3_cf_intrVec_11 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  REG__3_cf_brIdx = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  REG__3_cf_crossPageIPFFix = _RAND_121[0:0];
  _RAND_122 = {2{`RANDOM}};
  REG__3_cf_runahead_checkpoint_id = _RAND_122[63:0];
  _RAND_123 = {1{`RANDOM}};
  REG__3_ctrl_src1Type = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  REG__3_ctrl_src2Type = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  REG__3_ctrl_fuType = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  REG__3_ctrl_fuOpType = _RAND_126[6:0];
  _RAND_127 = {1{`RANDOM}};
  REG__3_ctrl_rfSrc1 = _RAND_127[4:0];
  _RAND_128 = {1{`RANDOM}};
  REG__3_ctrl_rfSrc2 = _RAND_128[4:0];
  _RAND_129 = {1{`RANDOM}};
  REG__3_ctrl_rfWen = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  REG__3_ctrl_rfDest = _RAND_130[4:0];
  _RAND_131 = {1{`RANDOM}};
  REG__3_ctrl_vtag = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  REG__3_ctrl_vec_addr = _RAND_132[4:0];
  _RAND_133 = {1{`RANDOM}};
  REG__3_ctrl_length_k = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  REG__3_ctrl_algorithm = _RAND_134[1:0];
  _RAND_135 = {2{`RANDOM}};
  REG__3_data_imm = _RAND_135[63:0];
  _RAND_136 = {1{`RANDOM}};
  REG_1 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  REG_2 = _RAND_137[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  output        io_out_mem_resp_ready,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_out_coh_req_ready,
  output        io_out_coh_req_valid,
  output [31:0] io_out_coh_req_bits_addr,
  output [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_ready,
  input         io_out_coh_resp_valid,
  input  [3:0]  io_out_coh_resp_bits_cmd,
  input  [63:0] io_out_coh_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[Coherence.scala 46:24]
  wire  _T_1 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_14 = ~inflight; // @[Coherence.scala 52:42]
  wire  _T_20 = ~inflight & _T_4; // @[Coherence.scala 52:52]
  reg [31:0] reqLatch_addr; // @[Reg.scala 15:16]
  reg [3:0] reqLatch_cmd; // @[Reg.scala 15:16]
  reg [63:0] reqLatch_wdata; // @[Reg.scala 15:16]
  wire  _T_23 = io_in_req_valid & _T_14; // @[Coherence.scala 65:43]
  wire  _GEN_5 = _T_4 & _T_23; // @[Coherence.scala 63:24 67:39 68:26]
  wire  _GEN_6 = _T_4 & (io_out_coh_req_ready & _T_14); // @[Coherence.scala 62:17 67:39 69:19]
  wire  _GEN_7 = io_in_req_bits_cmd[0] & (io_in_req_valid & _T_14); // @[Coherence.scala 61:24 64:61 65:26]
  wire  _T_36 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_43 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [2:0] _GEN_10 = _T_43 ? 3'h5 : state; // @[Coherence.scala 45:22 78:{48,56}]
  wire  _T_45 = io_out_coh_resp_ready & io_out_coh_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_46 = io_out_coh_resp_bits_cmd == 4'hc; // @[SimpleBus.scala 92:26]
  wire [2:0] _T_47 = _T_46 ? 3'h2 : 3'h3; // @[Coherence.scala 83:21]
  wire  _T_50 = io_in_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [2:0] _GEN_14 = io_in_resp_valid & _T_50 ? 3'h0 : state; // @[Coherence.scala 45:22 89:{60,68}]
  wire  _T_53 = io_out_mem_req_ready & io_out_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_53 ? 3'h4 : state; // @[Coherence.scala 45:22 94:{36,44}]
  wire  _T_55 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_56 = io_out_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [2:0] _GEN_16 = _T_55 & _T_56 ? 3'h0 : state; // @[Coherence.scala 96:101 45:22 96:93]
  wire [2:0] _GEN_17 = _T_55 ? 3'h0 : state; // @[Coherence.scala 45:22 97:{57,65}]
  wire [2:0] _GEN_18 = 3'h5 == state ? _GEN_17 : state; // @[Coherence.scala 74:18 45:22]
  wire [2:0] _GEN_19 = 3'h4 == state ? _GEN_16 : _GEN_18; // @[Coherence.scala 74:18]
  wire [63:0] _GEN_20 = 3'h3 == state ? reqLatch_wdata : io_in_req_bits_wdata; // @[Coherence.scala 74:18 59:23 92:27]
  wire [3:0] _GEN_22 = 3'h3 == state ? reqLatch_cmd : io_in_req_bits_cmd; // @[Coherence.scala 74:18 59:23 92:27]
  wire [31:0] _GEN_24 = 3'h3 == state ? reqLatch_addr : io_in_req_bits_addr; // @[Coherence.scala 74:18 59:23 92:27]
  wire  _GEN_25 = 3'h3 == state | _GEN_7; // @[Coherence.scala 74:18 93:28]
  wire [2:0] _GEN_26 = 3'h3 == state ? _GEN_15 : _GEN_19; // @[Coherence.scala 74:18]
  wire [63:0] _GEN_27 = 3'h2 == state ? io_out_coh_resp_bits_rdata : io_out_mem_resp_bits_rdata; // @[Coherence.scala 72:14 74:18 88:16]
  wire [3:0] _GEN_28 = 3'h2 == state ? io_out_coh_resp_bits_cmd : io_out_mem_resp_bits_cmd; // @[Coherence.scala 72:14 74:18 88:16]
  wire  _GEN_29 = 3'h2 == state ? io_out_coh_resp_valid : io_out_mem_resp_valid; // @[Coherence.scala 72:14 74:18 88:16]
  wire [63:0] _GEN_32 = 3'h2 == state ? io_in_req_bits_wdata : _GEN_20; // @[Coherence.scala 74:18 59:23]
  wire [3:0] _GEN_34 = 3'h2 == state ? io_in_req_bits_cmd : _GEN_22; // @[Coherence.scala 74:18 59:23]
  wire [31:0] _GEN_36 = 3'h2 == state ? io_in_req_bits_addr : _GEN_24; // @[Coherence.scala 74:18 59:23]
  wire  _GEN_37 = 3'h2 == state ? _GEN_7 : _GEN_25; // @[Coherence.scala 74:18]
  wire [63:0] _GEN_39 = 3'h1 == state ? io_out_mem_resp_bits_rdata : _GEN_27; // @[Coherence.scala 72:14 74:18]
  wire [3:0] _GEN_40 = 3'h1 == state ? io_out_mem_resp_bits_cmd : _GEN_28; // @[Coherence.scala 72:14 74:18]
  wire  _GEN_41 = 3'h1 == state ? io_out_mem_resp_valid : _GEN_29; // @[Coherence.scala 72:14 74:18]
  wire [63:0] _GEN_43 = 3'h1 == state ? io_in_req_bits_wdata : _GEN_32; // @[Coherence.scala 74:18 59:23]
  wire [3:0] _GEN_45 = 3'h1 == state ? io_in_req_bits_cmd : _GEN_34; // @[Coherence.scala 74:18 59:23]
  wire [31:0] _GEN_47 = 3'h1 == state ? io_in_req_bits_addr : _GEN_36; // @[Coherence.scala 74:18 59:23]
  wire  _GEN_48 = 3'h1 == state ? _GEN_7 : _GEN_37; // @[Coherence.scala 74:18]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? io_out_mem_req_ready & _T_14 : _GEN_6; // @[Coherence.scala 64:61 66:19]
  assign io_in_resp_valid = 3'h0 == state ? io_out_mem_resp_valid : _GEN_41; // @[Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_cmd = 3'h0 == state ? io_out_mem_resp_bits_cmd : _GEN_40; // @[Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_rdata = 3'h0 == state ? io_out_mem_resp_bits_rdata : _GEN_39; // @[Coherence.scala 72:14 74:18]
  assign io_out_mem_req_valid = 3'h0 == state ? _GEN_7 : _GEN_48; // @[Coherence.scala 74:18]
  assign io_out_mem_req_bits_addr = 3'h0 == state ? io_in_req_bits_addr : _GEN_47; // @[Coherence.scala 74:18 59:23]
  assign io_out_mem_req_bits_cmd = 3'h0 == state ? io_in_req_bits_cmd : _GEN_45; // @[Coherence.scala 74:18 59:23]
  assign io_out_mem_req_bits_wdata = 3'h0 == state ? io_in_req_bits_wdata : _GEN_43; // @[Coherence.scala 74:18 59:23]
  assign io_out_mem_resp_ready = 1'h1; // @[Coherence.scala 72:14]
  assign io_out_coh_req_valid = io_in_req_bits_cmd[0] ? 1'h0 : _GEN_5; // @[Coherence.scala 63:24 64:61]
  assign io_out_coh_req_bits_addr = io_in_req_bits_addr; // @[Coherence.scala 54:16]
  assign io_out_coh_req_bits_wdata = io_in_req_bits_wdata; // @[Coherence.scala 54:16]
  assign io_out_coh_resp_ready = 1'h1; // @[Coherence.scala 56:18 74:18]
  always @(posedge clock) begin
    if (reset) begin // @[Coherence.scala 45:22]
      state <= 3'h0; // @[Coherence.scala 45:22]
    end else if (3'h0 == state) begin // @[Coherence.scala 74:18]
      if (_T_36) begin // @[Coherence.scala 76:29]
        if (_T_4) begin // @[Coherence.scala 77:38]
          state <= 3'h1; // @[Coherence.scala 77:46]
        end else begin
          state <= _GEN_10;
        end
      end
    end else if (3'h1 == state) begin // @[Coherence.scala 74:18]
      if (_T_45) begin // @[Coherence.scala 82:37]
        state <= _T_47; // @[Coherence.scala 83:15]
      end
    end else if (3'h2 == state) begin // @[Coherence.scala 74:18]
      state <= _GEN_14;
    end else begin
      state <= _GEN_26;
    end
    if (_T_20) begin // @[Reg.scala 16:19]
      reqLatch_addr <= io_in_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (_T_20) begin // @[Reg.scala 16:19]
      reqLatch_cmd <= io_in_req_bits_cmd; // @[Reg.scala 16:23]
    end
    if (_T_20) begin // @[Reg.scala 16:19]
      reqLatch_wdata <= io_in_req_bits_wdata; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_req_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Coherence.scala:49 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Coherence.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_req_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Coherence.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqLatch_cmd = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  reqLatch_wdata = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI42SimpleBusConverter(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  input  [31:0] io_in_awaddr,
  input  [17:0] io_in_awid,
  input  [7:0]  io_in_awlen,
  input  [2:0]  io_in_awsize,
  output        io_in_wready,
  input         io_in_wvalid,
  input  [63:0] io_in_wdata,
  input  [7:0]  io_in_wstrb,
  input         io_in_wlast,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input  [17:0] io_in_arid,
  input  [7:0]  io_in_arlen,
  input  [2:0]  io_in_arsize,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata,
  output        io_in_rlast,
  output [17:0] io_in_rid,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] inflight_id_reg; // @[ToAXI4.scala 38:32]
  reg [1:0] inflight_type; // @[ToAXI4.scala 40:30]
  wire  _T = inflight_type == 2'h0; // @[ToAXI4.scala 50:19]
  wire  _T_1 = ~_T; // @[ToAXI4.scala 53:5]
  wire  _T_2 = ~_T_1; // @[ToAXI4.scala 64:9]
  wire  _T_3 = ~_T_1 & io_in_arvalid; // @[ToAXI4.scala 64:23]
  wire [1:0] _T_5 = io_in_arlen == 8'h0 ? 2'h0 : 2'h2; // @[ToAXI4.scala 67:19]
  wire  _T_6 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [17:0] _GEN_0 = _T_6 ? io_in_arid : inflight_id_reg; // @[ToAXI4.scala 42:21 74:25 38:32]
  wire [1:0] _GEN_1 = _T_6 ? 2'h1 : inflight_type; // @[ToAXI4.scala 43:19 74:25 40:30]
  wire [31:0] _GEN_2 = ~_T_1 & io_in_arvalid ? io_in_araddr : 32'h0; // @[ToAXI4.scala 64:40 66:14 59:7]
  wire [3:0] _GEN_3 = ~_T_1 & io_in_arvalid ? {{2'd0}, _T_5} : 4'h0; // @[ToAXI4.scala 64:40 67:13 59:7]
  wire [2:0] _GEN_4 = ~_T_1 & io_in_arvalid ? io_in_arsize : 3'h0; // @[ToAXI4.scala 64:40 69:14 59:7]
  wire [17:0] _GEN_7 = ~_T_1 & io_in_arvalid ? _GEN_0 : inflight_id_reg; // @[ToAXI4.scala 38:32 64:40]
  wire [1:0] _GEN_8 = ~_T_1 & io_in_arvalid ? _GEN_1 : inflight_type; // @[ToAXI4.scala 40:30 64:40]
  wire  _T_7 = inflight_type == 2'h1; // @[ToAXI4.scala 50:19]
  wire  _T_9 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_10 = io_in_rready & io_in_rvalid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_9 = _T_10 & _T_9 ? 2'h0 : _GEN_8; // @[ToAXI4.scala 46:19 88:42]
  wire [17:0] _GEN_10 = _T_10 & _T_9 ? 18'h0 : _GEN_7; // @[ToAXI4.scala 47:21 88:42]
  wire [1:0] _GEN_15 = _T_7 & io_out_resp_valid ? _GEN_9 : _GEN_8; // @[ToAXI4.scala 79:46]
  wire [17:0] _GEN_16 = _T_7 & io_out_resp_valid ? _GEN_10 : _GEN_7; // @[ToAXI4.scala 79:46]
  reg [31:0] aw_reg_addr; // @[ToAXI4.scala 94:19]
  reg [7:0] aw_reg_len; // @[ToAXI4.scala 94:19]
  reg [2:0] aw_reg_size; // @[ToAXI4.scala 94:19]
  reg  bresp_en; // @[ToAXI4.scala 95:25]
  wire  _T_17 = ~io_in_arvalid; // @[ToAXI4.scala 97:42]
  wire  _T_19 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_20 = inflight_type == 2'h2; // @[ToAXI4.scala 50:19]
  wire  _T_21 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_24 = io_in_wlast ? 3'h7 : 3'h3; // @[ToAXI4.scala 108:10]
  wire [2:0] _T_25 = aw_reg_len == 8'h0 ? 3'h1 : _T_24; // @[ToAXI4.scala 107:19]
  wire  _GEN_31 = io_in_wlast | bresp_en; // @[ToAXI4.scala 115:19 116:16 95:25]
  wire  _T_26 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  wire  _T_57 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_81 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  assign io_in_awready = _T_2 & _T_17; // @[ToAXI4.scala 132:33]
  assign io_in_wready = _T_20 & io_out_req_ready; // @[ToAXI4.scala 133:38]
  assign io_in_bvalid = bresp_en & io_out_resp_valid; // @[ToAXI4.scala 134:27]
  assign io_in_arready = _T_2 & io_out_req_ready; // @[ToAXI4.scala 129:33]
  assign io_in_rvalid = _T_7 & io_out_resp_valid; // @[ToAXI4.scala 130:36]
  assign io_in_rdata = _T_7 & io_out_resp_valid ? io_out_resp_bits_rdata : 64'h0; // @[ToAXI4.scala 79:46 81:12 60:5]
  assign io_in_rlast = _T_7 & io_out_resp_valid & _T_9; // @[ToAXI4.scala 79:46 85:12 60:5]
  assign io_in_rid = _T_7 & io_out_resp_valid ? inflight_id_reg : 18'h0; // @[ToAXI4.scala 79:46 82:10 60:5]
  assign io_out_req_valid = _T_3 | _T_20 & io_in_wvalid; // @[ToAXI4.scala 127:52]
  assign io_out_req_bits_addr = _T_20 & _T_21 ? aw_reg_addr : _GEN_2; // @[ToAXI4.scala 105:45 109:14]
  assign io_out_req_bits_size = _T_20 & _T_21 ? aw_reg_size : _GEN_4; // @[ToAXI4.scala 105:45 110:14]
  assign io_out_req_bits_cmd = _T_20 & _T_21 ? {{1'd0}, _T_25} : _GEN_3; // @[ToAXI4.scala 105:45 107:13]
  assign io_out_req_bits_wmask = _T_20 & _T_21 ? io_in_wstrb : 8'h0; // @[ToAXI4.scala 105:45 111:15]
  assign io_out_req_bits_wdata = _T_20 & _T_21 ? io_in_wdata : 64'h0; // @[ToAXI4.scala 105:45 112:15]
  assign io_out_resp_ready = _T_2 | _T_7 & io_in_rready | _T_20 & io_in_bready; // @[ToAXI4.scala 128:73]
  always @(posedge clock) begin
    if (reset) begin // @[ToAXI4.scala 38:32]
      inflight_id_reg <= 18'h0; // @[ToAXI4.scala 38:32]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      inflight_id_reg <= 18'h0; // @[ToAXI4.scala 47:21]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      if (_T_19) begin // @[ToAXI4.scala 100:24]
        inflight_id_reg <= io_in_awid; // @[ToAXI4.scala 42:21]
      end else begin
        inflight_id_reg <= _GEN_16;
      end
    end else begin
      inflight_id_reg <= _GEN_16;
    end
    if (reset) begin // @[ToAXI4.scala 40:30]
      inflight_type <= 2'h0; // @[ToAXI4.scala 40:30]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      inflight_type <= 2'h0; // @[ToAXI4.scala 46:19]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      if (_T_19) begin // @[ToAXI4.scala 100:24]
        inflight_type <= 2'h2; // @[ToAXI4.scala 43:19]
      end else begin
        inflight_type <= _GEN_15;
      end
    end else begin
      inflight_type <= _GEN_15;
    end
    if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_addr <= io_in_awaddr; // @[ToAXI4.scala 98:12]
    end
    if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_len <= io_in_awlen; // @[ToAXI4.scala 98:12]
    end
    if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_size <= io_in_awsize; // @[ToAXI4.scala 98:12]
    end
    if (reset) begin // @[ToAXI4.scala 95:25]
      bresp_en <= 1'h0; // @[ToAXI4.scala 95:25]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      bresp_en <= 1'h0; // @[ToAXI4.scala 121:14]
    end else if (_T_20 & _T_21) begin // @[ToAXI4.scala 105:45]
      bresp_en <= _GEN_31;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_57 & ~(_T_6 & _T_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:137 when (axi.ar.fire()) { assert(mem.req.fire() && !isInflight()); }\n"
            ); // @[ToAXI4.scala 137:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_57 & ~(_T_6 & _T_2 | reset)) begin
          $fatal; // @[ToAXI4.scala 137:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & ~(_T_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:138 when (axi.aw.fire()) { assert(!isInflight()); }\n"); // @[ToAXI4.scala 138:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_19 & ~(_T_2 | reset)) begin
          $fatal; // @[ToAXI4.scala 138:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & ~(_T_6 & _T_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:139 when (axi.w.fire()) { assert(mem.req .fire() && isState(axi_write)); }\n"
            ); // @[ToAXI4.scala 139:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_21 & ~(_T_6 & _T_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 139:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_26 & ~(_T_81 & _T_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:140 when (axi.b.fire()) { assert(mem.resp.fire() && isState(axi_write)); }\n"
            ); // @[ToAXI4.scala 140:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_26 & ~(_T_81 & _T_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 140:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(_T_81 & _T_7 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:141 when (axi.r.fire()) { assert(mem.resp.fire() && isState(axi_read)); }\n"
            ); // @[ToAXI4.scala 141:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10 & ~(_T_81 & _T_7 | reset)) begin
          $fatal; // @[ToAXI4.scala 141:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inflight_id_reg = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  inflight_type = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  aw_reg_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  aw_reg_len = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  aw_reg_size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  bresp_en = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Prefetcher(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  getNewReq; // @[Prefetcher.scala 37:26]
  reg [31:0] prefetchReq_addr; // @[Prefetcher.scala 38:28]
  reg [2:0] prefetchReq_size; // @[Prefetcher.scala 38:28]
  reg [7:0] prefetchReq_wmask; // @[Prefetcher.scala 38:28]
  reg [63:0] prefetchReq_wdata; // @[Prefetcher.scala 38:28]
  reg [63:0] lastReqAddr; // @[Prefetcher.scala 44:28]
  wire  _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_9 = {{32'd0}, io_in_bits_addr}; // @[Prefetcher.scala 50:30]
  wire [63:0] _T_4 = _GEN_9 & 64'hffffffffffffffc0; // @[Prefetcher.scala 50:30]
  wire [63:0] _T_5 = lastReqAddr & 64'hffffffffffffffc0; // @[Prefetcher.scala 50:59]
  wire  neqAddr = _T_4 != _T_5; // @[Prefetcher.scala 50:42]
  wire  _T_8 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _T_14 = prefetchReq_addr ^ 32'h30000000; // @[NutCore.scala 87:11]
  wire  _T_16 = _T_14[31:28] == 4'h0; // @[NutCore.scala 87:44]
  wire [31:0] _T_17 = prefetchReq_addr ^ 32'h40600000; // @[NutCore.scala 87:11]
  wire  _T_19 = _T_17[31:24] == 8'h0; // @[NutCore.scala 87:44]
  wire  _T_20 = _T_16 | _T_19; // @[NutCore.scala 88:15]
  assign io_in_ready = ~getNewReq & (~io_in_valid | _T_8); // @[Prefetcher.scala 52:21 55:17 60:17]
  assign io_out_valid = ~getNewReq ? io_in_valid : ~_T_20; // @[Prefetcher.scala 52:21 54:18 59:18]
  assign io_out_bits_addr = ~getNewReq ? io_in_bits_addr : prefetchReq_addr; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_size = ~getNewReq ? io_in_bits_size : prefetchReq_size; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_cmd = ~getNewReq ? io_in_bits_cmd : 4'h4; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_wmask = ~getNewReq ? io_in_bits_wmask : prefetchReq_wmask; // @[Prefetcher.scala 52:21 53:17 58:17]
  assign io_out_bits_wdata = ~getNewReq ? io_in_bits_wdata : prefetchReq_wdata; // @[Prefetcher.scala 52:21 53:17 58:17]
  always @(posedge clock) begin
    if (reset) begin // @[Prefetcher.scala 37:26]
      getNewReq <= 1'h0; // @[Prefetcher.scala 37:26]
    end else if (~getNewReq) begin // @[Prefetcher.scala 52:21]
      getNewReq <= _T_2 & io_in_bits_cmd[1] & neqAddr; // @[Prefetcher.scala 56:15]
    end else begin
      getNewReq <= ~(_T_8 | _T_20); // @[Prefetcher.scala 61:15]
    end
    prefetchReq_addr <= io_in_bits_addr + 32'h40; // @[Prefetcher.scala 40:39]
    prefetchReq_size <= io_in_bits_size; // @[Prefetcher.scala 38:28]
    prefetchReq_wmask <= io_in_bits_wmask; // @[Prefetcher.scala 38:28]
    prefetchReq_wdata <= io_in_bits_wdata; // @[Prefetcher.scala 38:28]
    if (reset) begin // @[Prefetcher.scala 44:28]
      lastReqAddr <= 64'h0; // @[Prefetcher.scala 44:28]
    end else if (_T_2) begin // @[Prefetcher.scala 45:23]
      lastReqAddr <= {{32'd0}, io_in_bits_addr}; // @[Prefetcher.scala 46:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  getNewReq = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  prefetchReq_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  prefetchReq_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  prefetchReq_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  prefetchReq_wdata = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  lastReqAddr = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheStage1_2(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [8:0]  io_metaReadBus_req_bits_setIdx,
  input  [16:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [16:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [16:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [16:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_16 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_16) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 147:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 146:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 145:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 145:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 145:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 145:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[14:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 141:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[14:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module CacheStage2_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [16:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_dirty,
  output [16:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_dirty,
  output [16:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_dirty,
  output [16:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [16:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [16:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [16:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [16:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [8:0]  io_metaWriteBus_req_bits_setIdx,
  input  [16:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [11:0] io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 176:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 176:31]
  wire [16:0] addr_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 176:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 178:64]
  reg  isForwardMetaReg; // @[Cache.scala 179:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 180:24 179:33 180:43]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 181:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 181:22]
  reg [16:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 15:16 16:{19,23}]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 15:16 16:{19,23}]
  wire [16:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 15:16 16:{19,23}]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 185:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 187:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 187:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 187:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 187:61]
  wire [16:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 | io_metaReadResp_0_valid; // @[Cache.scala 189:22]
  wire [16:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 | io_metaReadResp_1_valid; // @[Cache.scala 189:22]
  wire [16:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 | io_metaReadResp_2_valid; // @[Cache.scala 189:22]
  wire [16:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 | io_metaReadResp_3_valid; // @[Cache.scala 189:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 192:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 192:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  _T_39 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _T_42 = {_T_39,REG[63:1]}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 193:42]
  wire  _T_45 = ~metaWay_0_valid; // @[Cache.scala 195:45]
  wire  _T_46 = ~metaWay_1_valid; // @[Cache.scala 195:45]
  wire  _T_47 = ~metaWay_2_valid; // @[Cache.scala 195:45]
  wire  _T_48 = ~metaWay_3_valid; // @[Cache.scala 195:45]
  wire [3:0] invalidVec = {_T_48,_T_47,_T_46,_T_45}; // @[Cache.scala 195:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 196:34]
  wire [1:0] _T_52 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 199:8]
  wire [2:0] _T_53 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_52}; // @[Cache.scala 198:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_53}; // @[Cache.scala 197:33]
  wire [3:0] _T_54 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 202:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  wire [1:0] _T_59 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_61 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_63 = _T_59 + _T_61; // @[Bitwise.scala 47:55]
  wire  _T_65 = _T_63 > 3'h1; // @[Cache.scala 203:26]
  wire [31:0] _T_172 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 87:11]
  wire  _T_174 = _T_172[31:28] == 4'h0; // @[NutCore.scala 87:44]
  wire [31:0] _T_175 = io_in_bits_req_addr ^ 32'h40600000; // @[NutCore.scala 87:11]
  wire  _T_177 = _T_175[31:24] == 8'h0; // @[NutCore.scala 87:44]
  wire [11:0] _T_187 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_189 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_187; // @[Cache.scala 219:13]
  wire  isForwardData = io_in_valid & _T_189; // @[Cache.scala 218:35]
  reg  isForwardDataReg; // @[Cache.scala 221:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 222:24 221:33 222:43]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_196 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_196; // @[Cache.scala 230:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 229:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 228:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 228:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 228:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 228:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 189:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 189:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 215:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 215:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 213:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_54; // @[Cache.scala 202:20]
  assign io_out_bits_mmio = _T_174 | _T_177; // @[NutCore.scala 88:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 225:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 226:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 226:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 179:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 179:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 181:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 181:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[Reg.scala 16:23]
    end
    if (isForwardMeta) begin // @[Reg.scala 16:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_42;
    end
    if (reset) begin // @[Cache.scala 221:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 221:33]
    end else if (_T_12) begin // @[Cache.scala 223:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 223:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 16:23]
    end
    if (isForwardData) begin // @[Reg.scala 16:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:210 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 210:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_65) | reset)) begin
          $fatal; // @[Cache.scala 210:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  REG = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_10(
  input         io_in_0_valid,
  input  [8:0]  io_in_0_bits_setIdx,
  input  [16:0] io_in_0_bits_data_tag,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [8:0]  io_in_1_bits_setIdx,
  input  [16:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [8:0]  io_out_bits_setIdx,
  output [16:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid | io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module Arbiter_11(
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 126:27 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module CacheStage3_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [16:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_dirty,
  input  [16:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_dirty,
  input  [16:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_dirty,
  input  [16:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [11:0] io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [8:0]  io_metaWriteBus_req_bits_setIdx,
  output [16:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  output        io_cohResp_valid,
  output        io_dataReadRespToL1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 256:28]
  wire [8:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 256:28]
  wire [16:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 256:28]
  wire [8:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 256:28]
  wire [16:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 256:28]
  wire [8:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 256:28]
  wire [16:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 256:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 256:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 256:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 257:28]
  wire [11:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 257:28]
  wire [11:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 257:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 257:28]
  wire [11:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 257:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 257:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 257:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 260:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 260:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 261:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 262:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 263:26]
  wire  _T_6 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_6; // @[Cache.scala 264:39]
  wire  _T_7 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_7; // @[Cache.scala 265:26]
  wire  meta_dirty = io_in_bits_waymask[0] & io_in_bits_metas_0_dirty | io_in_bits_waymask[1] & io_in_bits_metas_1_dirty
     | io_in_bits_waymask[2] & io_in_bits_metas_2_dirty | io_in_bits_waymask[3] & io_in_bits_metas_3_dirty; // @[Mux.scala 27:72]
  wire [16:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 17'h0; // @[Mux.scala 27:72]
  wire [16:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [16:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [16:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 275:49]
  wire [63:0] _T_43 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_43 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_48 | _T_46; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_49; // @[Cache.scala 277:21]
  wire [7:0] _T_62 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_64 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_66 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_77 = {_T_76,_T_74,_T_72,_T_70,_T_68,_T_66,_T_64,_T_62}; // @[Cat.scala 30:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_77 : 64'h0; // @[Cache.scala 278:21]
  reg [2:0] value; // @[Counter.scala 60:40]
  wire  _T_79 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 281:34]
  wire  _T_80 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_81 = io_in_bits_req_cmd == 4'h3 | _T_80; // @[Cache.scala 281:62]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_0 = io_out_valid & (io_in_bits_req_cmd == 4'h3 | _T_80) ? _value_T_1 : value; // @[Cache.scala 281:85 Counter.scala 76:15 60:40]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 285:22]
  wire [63:0] _T_84 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_85 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_86 = dataRead & _T_85; // @[BitUtils.scala 32:36]
  wire [2:0] _T_91 = _T_81 ? value : addr_wordIndex; // @[Cache.scala 288:51]
  wire  metaHitWriteBus_req_valid = hitWrite & ~meta_dirty; // @[Cache.scala 291:22]
  reg [3:0] state; // @[Cache.scala 296:22]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 306:23]
  wire  _T_103 = state == 4'h3; // @[Cache.scala 308:39]
  wire  _T_104 = state == 4'h8; // @[Cache.scala 308:66]
  wire [2:0] _T_109 = _T_104 ? value_1 : value_2; // @[Cache.scala 309:33]
  wire  _T_111 = state2 == 2'h1; // @[Cache.scala 310:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_116 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_117 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_118 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_119 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_120 = _T_116 | _T_117; // @[Mux.scala 27:72]
  wire [63:0] _T_121 = _T_120 | _T_118; // @[Mux.scala 27:72]
  wire [63:0] _T_122 = _T_121 | _T_119; // @[Mux.scala 27:72]
  wire  _T_124 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_127 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_8 = _T_127 | io_cohResp_valid | hitReadBurst ? 2'h0 : state2; // @[Cache.scala 316:{100,109} 306:23]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_133 = state == 4'h1; // @[Cache.scala 324:23]
  wire [2:0] _T_135 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 325:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_135; // @[Cache.scala 324:16]
  wire  _T_141 = state2 == 2'h2; // @[Cache.scala 331:89]
  reg  afterFirstRead; // @[Cache.scala 338:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = io_out_valid | alreadyOutFire; // @[Reg.scala 28:19 27:20 28:23]
  wire  _T_147 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_149 = state == 4'h2; // @[Cache.scala 340:70]
  wire  readingFirst = ~afterFirstRead & _T_147 & state == 4'h2; // @[Cache.scala 340:60]
  wire  _T_152 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 342:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_153 = state == 4'h0; // @[Cache.scala 345:31]
  wire  _T_157 = _T_104 & _T_141; // @[Cache.scala 346:46]
  wire  _T_161 = _T_104 & io_cohResp_valid; // @[Cache.scala 348:49]
  reg [2:0] value_3; // @[Counter.scala 60:40]
  wire  wrap_wrap = value_3 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_1 = value_3 + 3'h1; // @[Counter.scala 76:24]
  wire  releaseLast = _T_161 & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  respToL1Fire = hitReadBurst & _T_141; // @[Cache.scala 352:51]
  wire  _T_172 = _T_153 | _T_157; // @[Cache.scala 353:48]
  wire  _T_173 = (_T_153 | _T_157) & hitReadBurst; // @[Cache.scala 353:96]
  reg [2:0] value_4; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = value_4 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_3 = value_4 + 3'h1; // @[Counter.scala 76:24]
  wire  respToL1Last = _T_173 & wrap_wrap_1; // @[Counter.scala 118:{17,24}]
  wire [3:0] _T_177 = hit ? 4'h8 : 4'h0; // @[Cache.scala 362:23]
  wire [2:0] _value_T_4 = addr_wordIndex + 3'h1; // @[Cache.scala 367:93]
  wire [2:0] _value_T_5 = addr_wordIndex == 3'h7 ? 3'h0 : _value_T_4; // @[Cache.scala 367:33]
  wire [3:0] _T_184 = meta_dirty ? 4'h3 : 4'h1; // @[Cache.scala 369:42]
  wire [3:0] _T_185 = mmio ? 4'h5 : _T_184; // @[Cache.scala 369:21]
  wire [3:0] _GEN_20 = miss | mmio ? _T_185 : state; // @[Cache.scala 368:49 369:15 296:22]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid | respToL1Fire ? _value_T_7 : value_1; // @[Cache.scala 377:48 Counter.scala 76:15 60:40]
  wire  _T_196 = respToL1Fire & respToL1Last; // @[Cache.scala 378:71]
  wire [3:0] _GEN_28 = probe & io_cohResp_valid & releaseLast | respToL1Fire & respToL1Last ? 4'h0 : state; // @[Cache.scala 296:22 378:{88,96}]
  wire [3:0] _GEN_29 = _T_127 ? 4'h2 : state; // @[Cache.scala 381:50 382:13 296:22]
  wire [2:0] _GEN_30 = _T_127 ? addr_wordIndex : value_1; // @[Cache.scala 381:50 383:25 Counter.scala 60:40]
  wire [2:0] _GEN_31 = _T_79 ? 3'h0 : _GEN_0; // @[Cache.scala 390:{52,75}]
  wire  _T_203 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_203 ? 4'h7 : state; // @[Cache.scala 296:22 391:{46,54}]
  wire  _GEN_33 = _T_147 | afterFirstRead; // @[Cache.scala 387:33 388:24 338:31]
  wire [2:0] _GEN_34 = _T_147 ? _value_T_7 : value_1; // @[Cache.scala 387:33 Counter.scala 76:15 60:40]
  wire [2:0] _GEN_35 = _T_147 ? _GEN_31 : _GEN_0; // @[Cache.scala 387:33]
  wire [3:0] _GEN_36 = _T_147 ? _GEN_32 : state; // @[Cache.scala 296:22 387:33]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_127 ? _value_T_11 : value_2; // @[Cache.scala 396:32 Counter.scala 76:15 60:40]
  wire  _T_206 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_206 & _T_127 ? 4'h4 : state; // @[Cache.scala 296:22 397:{65,73}]
  wire [3:0] _GEN_39 = _T_147 ? 4'h1 : state; // @[Cache.scala 296:22 400:{53,61}]
  wire [3:0] _GEN_40 = _GEN_12 ? 4'h0 : state; // @[Cache.scala 296:22 401:{76,84}]
  wire [3:0] _GEN_41 = 4'h7 == state ? _GEN_40 : state; // @[Cache.scala 355:18 296:22]
  wire [3:0] _GEN_42 = 4'h4 == state ? _GEN_39 : _GEN_41; // @[Cache.scala 355:18]
  wire [2:0] _GEN_43 = 4'h3 == state ? _GEN_37 : value_2; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [3:0] _GEN_44 = 4'h3 == state ? _GEN_38 : _GEN_42; // @[Cache.scala 355:18]
  wire  _GEN_45 = 4'h2 == state ? _GEN_33 : afterFirstRead; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_46 = 4'h2 == state ? _GEN_34 : value_1; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [2:0] _GEN_47 = 4'h2 == state ? _GEN_35 : _GEN_0; // @[Cache.scala 355:18]
  wire [3:0] _GEN_48 = 4'h2 == state ? _GEN_36 : _GEN_44; // @[Cache.scala 355:18]
  wire [2:0] _GEN_49 = 4'h2 == state ? value_2 : _GEN_43; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [3:0] _GEN_50 = 4'h1 == state ? _GEN_29 : _GEN_48; // @[Cache.scala 355:18]
  wire [2:0] _GEN_51 = 4'h1 == state ? _GEN_30 : _GEN_46; // @[Cache.scala 355:18]
  wire  _GEN_52 = 4'h1 == state ? afterFirstRead : _GEN_45; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_53 = 4'h1 == state ? _GEN_0 : _GEN_47; // @[Cache.scala 355:18]
  wire [2:0] _GEN_54 = 4'h1 == state ? value_2 : _GEN_49; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [2:0] _GEN_55 = 4'h8 == state ? _GEN_27 : _GEN_51; // @[Cache.scala 355:18]
  wire [3:0] _GEN_56 = 4'h8 == state ? _GEN_28 : _GEN_50; // @[Cache.scala 355:18]
  wire  _GEN_57 = 4'h8 == state ? afterFirstRead : _GEN_52; // @[Cache.scala 355:18 338:31]
  wire [2:0] _GEN_58 = 4'h8 == state ? _GEN_0 : _GEN_53; // @[Cache.scala 355:18]
  wire [2:0] _GEN_59 = 4'h8 == state ? value_2 : _GEN_54; // @[Cache.scala 355:18 Counter.scala 60:40]
  wire [63:0] _T_215 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 404:67]
  wire [63:0] _T_216 = io_in_bits_req_wdata & _T_215; // @[BitUtils.scala 32:13]
  wire [63:0] _T_217 = ~_T_215; // @[BitUtils.scala 32:38]
  wire [63:0] _T_218 = io_mem_resp_bits_rdata & _T_217; // @[BitUtils.scala 32:36]
  wire [63:0] dataRefill = _T_216 | _T_218; // @[BitUtils.scala 32:25]
  wire  dataRefillWriteBus_req_valid = _T_149 & _T_147; // @[Cache.scala 406:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_203; // @[Cache.scala 414:61]
  wire  _T_239 = dataRefillWriteBus_req_valid & _T_7; // @[Cache.scala 424:59]
  wire [2:0] _T_241 = _T_203 ? 3'h6 : 3'h2; // @[Cache.scala 427:29]
  wire [63:0] _T_245 = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 430:31]
  wire [2:0] _T_248 = respToL1Last ? 3'h6 : 3'h2; // @[Cache.scala 435:29]
  wire [63:0] _GEN_76 = hitReadBurst & _T_104 ? _T_122 : _T_245; // @[Cache.scala 432:54 434:25 437:25]
  wire [3:0] _GEN_77 = hitReadBurst & _T_104 ? {{1'd0}, _T_248} : io_in_bits_req_cmd; // @[Cache.scala 432:54 435:23 438:23]
  wire [63:0] _GEN_78 = _T_80 | _T_79 ? _T_245 : _GEN_76; // @[Cache.scala 428:75 430:25]
  wire  _T_254 = state == 4'h7; // @[Cache.scala 448:48]
  wire  _T_267 = io_in_bits_req_cmd[0] & (hit | ~hit & state == 4'h7) | _T_239 | _T_196 & _T_104; // @[Cache.scala 448:161]
  wire  _T_273 = io_in_bits_req_cmd[0] | mmio ? _T_254 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 449:45]
  wire  _T_275 = probe ? 1'h0 : hit | _T_273; // @[Cache.scala 449:8]
  wire  _T_276 = io_in_bits_req_cmd[1] ? _T_267 : _T_275; // @[Cache.scala 447:37]
  wire  _T_282 = miss ? _T_153 : _T_104 & releaseLast; // @[Cache.scala 456:53]
  wire  _T_291 = hit | io_in_bits_req_cmd[0] ? io_out_valid : _T_254 & _GEN_12; // @[Cache.scala 457:8]
  Arbiter_10 metaWriteArb ( // @[Cache.scala 256:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_11 dataWriteArb ( // @[Cache.scala 257:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_153 & ~hitReadBurst & ~miss & ~probe; // @[Cache.scala 460:79]
  assign io_out_valid = io_in_valid & _T_276; // @[Cache.scala 447:31]
  assign io_out_bits_cmd = dataRefillWriteBus_req_valid & _T_7 ? {{1'd0}, _T_241} : _GEN_77; // @[Cache.scala 424:81 427:23]
  assign io_out_bits_rdata = dataRefillWriteBus_req_valid & _T_7 ? dataRefill : _GEN_78; // @[Cache.scala 424:81 426:25]
  assign io_isFinish = probe ? io_cohResp_valid & _T_282 : _T_291; // @[Cache.scala 456:21]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 308:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_109}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 411:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 411:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 421:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 421:23]
  assign io_mem_req_valid = _T_133 | _T_103 & state2 == 2'h2; // @[Cache.scala 331:48]
  assign io_mem_req_bits_addr = _T_133 ? raddr : waddr; // @[Cache.scala 326:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_121 | _T_119; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 330:21]
  assign io_cohResp_valid = state == 4'h0 & probe | _T_157; // @[Cache.scala 345:53]
  assign io_dataReadRespToL1 = hitReadBurst & _T_172; // @[Cache.scala 461:39]
  assign metaWriteArb_io_in_0_valid = hitWrite & ~meta_dirty; // @[Cache.scala 291:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 290:29 SRAMTemplate.scala 38:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_203; // @[Cache.scala 414:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 260:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[SimpleBus.scala 74:22]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 413:32 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 285:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_91}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = _T_84 | _T_86; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 286:29 SRAMTemplate.scala 38:24]
  assign dataWriteArb_io_in_1_valid = _T_149 & _T_147; // @[Cache.scala 406:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = _T_216 | _T_218; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:32 SRAMTemplate.scala 38:24]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      value <= _GEN_0;
    end else if (4'h5 == state) begin // @[Cache.scala 355:18]
      value <= _GEN_0;
    end else if (4'h6 == state) begin // @[Cache.scala 355:18]
      value <= _GEN_0;
    end else begin
      value <= _GEN_58;
    end
    if (reset) begin // @[Cache.scala 296:22]
      state <= 4'h0; // @[Cache.scala 296:22]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      if (probe) begin // @[Cache.scala 360:20]
        if (io_cohResp_valid) begin // @[Cache.scala 361:34]
          state <= _T_177; // @[Cache.scala 362:17]
        end
      end else if (hitReadBurst) begin // @[Cache.scala 365:50]
        state <= 4'h8; // @[Cache.scala 366:15]
      end else begin
        state <= _GEN_20;
      end
    end else if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
        state <= _GEN_56;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      if (probe) begin // @[Cache.scala 360:20]
        if (io_cohResp_valid) begin // @[Cache.scala 361:34]
          value_1 <= addr_wordIndex; // @[Cache.scala 363:29]
        end
      end else if (hitReadBurst) begin // @[Cache.scala 365:50]
        value_1 <= _value_T_5; // @[Cache.scala 367:27]
      end
    end else if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
        value_1 <= _GEN_55;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
        if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 306:23]
      state2 <= 2'h0; // @[Cache.scala 306:23]
    end else if (2'h0 == state2) begin // @[Cache.scala 313:19]
      if (_T_124) begin // @[Cache.scala 314:53]
        state2 <= 2'h1; // @[Cache.scala 314:62]
      end
    end else if (2'h1 == state2) begin // @[Cache.scala 313:19]
      state2 <= 2'h2; // @[Cache.scala 315:35]
    end else if (2'h2 == state2) begin // @[Cache.scala 313:19]
      state2 <= _GEN_8;
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 16:23]
    end
    if (_T_111) begin // @[Reg.scala 16:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Cache.scala 338:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 338:31]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      afterFirstRead <= 1'h0; // @[Cache.scala 357:22]
    end else if (!(4'h5 == state)) begin // @[Cache.scala 355:18]
      if (!(4'h6 == state)) begin // @[Cache.scala 355:18]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (4'h0 == state) begin // @[Cache.scala 355:18]
      alreadyOutFire <= 1'h0; // @[Cache.scala 358:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_152) begin // @[Reg.scala 16:19]
      if (mmio) begin // @[Cache.scala 341:39]
        inRdataRegDemand <= 64'h0;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_3 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_161) begin // @[Counter.scala 118:17]
      value_3 <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_4 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_173) begin // @[Counter.scala 118:17]
      value_4 <= _wrap_value_T_3; // @[Counter.scala 76:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:267 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 267:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 267:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:463 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 463:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 463:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:464 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 464:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 464:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  value_3 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  value_4 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_5(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [8:0]  io_rreq_bits_setIdx,
  output [16:0] io_rresp_data_0_tag,
  output        io_rresp_data_0_valid,
  output        io_rresp_data_0_dirty,
  output [16:0] io_rresp_data_1_tag,
  output        io_rresp_data_1_valid,
  output        io_rresp_data_1_dirty,
  output [16:0] io_rresp_data_2_tag,
  output        io_rresp_data_2_valid,
  output        io_rresp_data_2_dirty,
  output [16:0] io_rresp_data_3_tag,
  output        io_rresp_data_3_valid,
  output        io_rresp_data_3_dirty,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [16:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  reg  REG; // @[SRAMTemplate.scala 80:30]
  reg [8:0] value; // @[Counter.scala 60:40]
  wire  wrap_wrap = value == 9'h1ff; // @[Counter.scala 72:24]
  wire [8:0] _wrap_value_T_1 = value + 9'h1; // @[Counter.scala 76:24]
  wire  wrap = REG & wrap_wrap; // @[Counter.scala 118:{17,24}]
  wire  _GEN_2 = wrap ? 1'h0 : REG; // @[SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  wire  _T = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 89:38]
  wire [8:0] setIdx = REG ? value : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [18:0] _T_1 = {io_wreq_bits_data_tag,1'h1,io_wreq_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = REG ? 4'hf : io_wreq_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [18:0] _WIRE_2 = array_RW0_rdata_0;
  wire [18:0] _WIRE_3 = array_RW0_rdata_1;
  wire [18:0] _WIRE_4 = array_RW0_rdata_2;
  wire [18:0] _WIRE_5 = array_RW0_rdata_3;
  array_2 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~REG & _T; // @[SRAMTemplate.scala 101:33]
  assign io_rresp_data_0_tag = _WIRE_2[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_valid = _WIRE_2[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_0_dirty = _WIRE_2[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_tag = _WIRE_3[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_valid = _WIRE_3[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_dirty = _WIRE_3[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_tag = _WIRE_4[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_valid = _WIRE_4[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_dirty = _WIRE_4[0]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_tag = _WIRE_5[18:2]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_valid = _WIRE_5[1]; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_dirty = _WIRE_5[0]; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = REG ? 19'h0 : _T_1; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | wen;
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[Counter.scala 60:40]
      value <= 9'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      value <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter_12(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [8:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [8:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter_4(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [8:0]  io_r0_req_bits_setIdx,
  output [16:0] io_r0_resp_data_0_tag,
  output        io_r0_resp_data_0_valid,
  output        io_r0_resp_data_0_dirty,
  output [16:0] io_r0_resp_data_1_tag,
  output        io_r0_resp_data_1_valid,
  output        io_r0_resp_data_1_dirty,
  output [16:0] io_r0_resp_data_2_tag,
  output        io_r0_resp_data_2_valid,
  output        io_r0_resp_data_2_dirty,
  output [16:0] io_r0_resp_data_3_tag,
  output        io_r0_resp_data_3_valid,
  output        io_r0_resp_data_3_dirty,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [16:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_wreq_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [16:0] r_0_tag; // @[Reg.scala 27:20]
  reg  r_0_valid; // @[Reg.scala 27:20]
  reg  r_0_dirty; // @[Reg.scala 27:20]
  reg [16:0] r_1_tag; // @[Reg.scala 27:20]
  reg  r_1_valid; // @[Reg.scala 27:20]
  reg  r_1_dirty; // @[Reg.scala 27:20]
  reg [16:0] r_2_tag; // @[Reg.scala 27:20]
  reg  r_2_valid; // @[Reg.scala 27:20]
  reg  r_2_dirty; // @[Reg.scala 27:20]
  reg [16:0] r_3_tag; // @[Reg.scala 27:20]
  reg  r_3_valid; // @[Reg.scala 27:20]
  reg  r_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_5 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(ram_io_rresp_data_0_tag),
    .io_rresp_data_0_valid(ram_io_rresp_data_0_valid),
    .io_rresp_data_0_dirty(ram_io_rresp_data_0_dirty),
    .io_rresp_data_1_tag(ram_io_rresp_data_1_tag),
    .io_rresp_data_1_valid(ram_io_rresp_data_1_valid),
    .io_rresp_data_1_dirty(ram_io_rresp_data_1_dirty),
    .io_rresp_data_2_tag(ram_io_rresp_data_2_tag),
    .io_rresp_data_2_valid(ram_io_rresp_data_2_valid),
    .io_rresp_data_2_dirty(ram_io_rresp_data_2_dirty),
    .io_rresp_data_3_tag(ram_io_rresp_data_3_tag),
    .io_rresp_data_3_valid(ram_io_rresp_data_3_valid),
    .io_rresp_data_3_dirty(ram_io_rresp_data_3_dirty),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(ram_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(ram_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_12 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_tag = REG ? ram_io_rresp_data_0_tag : r_0_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_valid = REG ? ram_io_rresp_data_0_valid : r_0_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_dirty = REG ? ram_io_rresp_data_0_dirty : r_0_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_tag = REG ? ram_io_rresp_data_1_tag : r_1_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_valid = REG ? ram_io_rresp_data_1_valid : r_1_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_dirty = REG ? ram_io_rresp_data_1_dirty : r_1_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_tag = REG ? ram_io_rresp_data_2_tag : r_2_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_valid = REG ? ram_io_rresp_data_2_valid : r_2_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_dirty = REG ? ram_io_rresp_data_2_dirty : r_2_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_tag = REG ? ram_io_rresp_data_3_tag : r_3_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_valid = REG ? ram_io_rresp_data_3_valid : r_3_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_dirty = REG ? ram_io_rresp_data_3_dirty : r_3_dirty; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_tag = io_wreq_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_dirty = io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_0_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_tag <= ram_io_rresp_data_0_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_valid <= ram_io_rresp_data_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_0_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_0_dirty <= ram_io_rresp_data_0_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_tag <= ram_io_rresp_data_1_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_valid <= ram_io_rresp_data_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_1_dirty <= ram_io_rresp_data_1_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_tag <= ram_io_rresp_data_2_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_valid <= ram_io_rresp_data_2_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_2_dirty <= ram_io_rresp_data_2_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_tag <= 17'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_tag <= ram_io_rresp_data_3_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_valid <= ram_io_rresp_data_3_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_3_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r_3_dirty <= ram_io_rresp_data_3_dirty; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_0_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  r_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1_tag = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  r_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_2_tag = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  r_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_3_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  r_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRAMTemplate_6(
  input         clock,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [11:0] io_rreq_bits_setIdx,
  output [63:0] io_rresp_data_0_data,
  output [63:0] io_rresp_data_1_data,
  output [63:0] io_rresp_data_2_data,
  output [63:0] io_rresp_data_3_data,
  input         io_wreq_valid,
  input  [11:0] io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
  wire [11:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  wire  realRen = io_rreq_valid & ~io_wreq_valid; // @[SRAMTemplate.scala 89:38]
  array_3 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~io_wreq_valid; // @[SRAMTemplate.scala 101:53]
  assign io_rresp_data_0_data = array_RW0_rdata_0; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_1_data = array_RW0_rdata_1; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_2_data = array_RW0_rdata_2; // @[SRAMTemplate.scala 98:78]
  assign io_rresp_data_3_data = array_RW0_rdata_3; // @[SRAMTemplate.scala 98:78]
  assign array_RW0_clk = clock; // @[SRAMTemplate.scala 95:14]
  assign array_RW0_wdata_0 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_1 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_2 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wdata_3 = io_wreq_bits_data_data; // @[SRAMTemplate.scala 92:22]
  assign array_RW0_wmask_0 = io_wreq_bits_waymask[0]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_1 = io_wreq_bits_waymask[1]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_2 = io_wreq_bits_waymask[2]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_wmask_3 = io_wreq_bits_waymask[3]; // @[SRAMTemplate.scala 95:51]
  assign array_RW0_en = realRen | io_wreq_valid;
  assign array_RW0_wmode = io_wreq_valid; // @[SRAMTemplate.scala 88:52]
  assign array_RW0_addr = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx;
endmodule
module Arbiter_13(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 126:27 128:19]
endmodule
module SRAMTemplateWithArbiter_5(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [11:0] io_r0_req_bits_setIdx,
  output [63:0] io_r0_resp_data_0_data,
  output [63:0] io_r0_resp_data_1_data,
  output [63:0] io_r0_resp_data_2_data,
  output [63:0] io_r0_resp_data_3_data,
  output        io_r1_req_ready,
  input         io_r1_req_valid,
  input  [11:0] io_r1_req_bits_setIdx,
  output [63:0] io_r1_resp_data_0_data,
  output [63:0] io_r1_resp_data_1_data,
  output [63:0] io_r1_resp_data_2_data,
  output [63:0] io_r1_resp_data_3_data,
  input         io_wreq_valid,
  input  [11:0] io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_wreq_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  REG; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r__0_data; // @[Reg.scala 27:20]
  reg [63:0] r__1_data; // @[Reg.scala 27:20]
  reg [63:0] r__2_data; // @[Reg.scala 27:20]
  reg [63:0] r__3_data; // @[Reg.scala 27:20]
  reg  REG_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] r_1_0_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_1_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_2_data; // @[Reg.scala 27:20]
  reg [63:0] r_1_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_6 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_data(ram_io_rresp_data_0_data),
    .io_rresp_data_1_data(ram_io_rresp_data_1_data),
    .io_rresp_data_2_data(ram_io_rresp_data_2_data),
    .io_rresp_data_3_data(ram_io_rresp_data_3_data),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(ram_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_13 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_data = REG ? ram_io_rresp_data_0_data : r__0_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_data = REG ? ram_io_rresp_data_1_data : r__1_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_data = REG ? ram_io_rresp_data_2_data : r__2_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_data = REG ? ram_io_rresp_data_3_data : r__3_data; // @[Hold.scala 23:48]
  assign io_r1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r1_resp_data_0_data = REG_1 ? ram_io_rresp_data_0_data : r_1_0_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_1_data = REG_1 ? ram_io_rresp_data_1_data : r_1_1_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_2_data = REG_1 ? ram_io_rresp_data_2_data : r_1_2_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_3_data = REG_1 ? ram_io_rresp_data_3_data : r_1_3_data; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_data = io_wreq_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
  always @(posedge clock) begin
    REG <= io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r__0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r__3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      r__3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
    REG_1 <= io_r1_req_ready & io_r1_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_1_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r_1_3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r__0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  r__1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  r__2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  r__3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r_1_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  r_1_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  r_1_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache_2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 482:18]
  wire  s1_io_in_valid; // @[Cache.scala 482:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 482:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 482:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 482:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 482:18]
  wire  s1_io_out_ready; // @[Cache.scala 482:18]
  wire  s1_io_out_valid; // @[Cache.scala 482:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 482:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 482:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 482:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 482:18]
  wire [8:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 482:18]
  wire [16:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 482:18]
  wire [16:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 482:18]
  wire [16:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 482:18]
  wire [16:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 482:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 482:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 482:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 482:18]
  wire [11:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 482:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 482:18]
  wire  s2_clock; // @[Cache.scala 483:18]
  wire  s2_reset; // @[Cache.scala 483:18]
  wire  s2_io_in_ready; // @[Cache.scala 483:18]
  wire  s2_io_in_valid; // @[Cache.scala 483:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 483:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 483:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 483:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 483:18]
  wire  s2_io_out_ready; // @[Cache.scala 483:18]
  wire  s2_io_out_valid; // @[Cache.scala 483:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 483:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 483:18]
  wire [16:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 483:18]
  wire [16:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 483:18]
  wire [16:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 483:18]
  wire [16:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 483:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 483:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 483:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 483:18]
  wire [16:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 483:18]
  wire [16:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 483:18]
  wire [16:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 483:18]
  wire [16:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 483:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 483:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 483:18]
  wire [8:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 483:18]
  wire [16:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 483:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 483:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 483:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 483:18]
  wire [11:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 483:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 483:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 483:18]
  wire  s3_clock; // @[Cache.scala 484:18]
  wire  s3_reset; // @[Cache.scala 484:18]
  wire  s3_io_in_ready; // @[Cache.scala 484:18]
  wire  s3_io_in_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 484:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 484:18]
  wire [16:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 484:18]
  wire [16:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 484:18]
  wire [16:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 484:18]
  wire [16:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 484:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 484:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 484:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 484:18]
  wire  s3_io_out_valid; // @[Cache.scala 484:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_isFinish; // @[Cache.scala 484:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 484:18]
  wire [11:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 484:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 484:18]
  wire [11:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 484:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 484:18]
  wire [8:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 484:18]
  wire [16:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 484:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 484:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 484:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 484:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 484:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 484:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 484:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 484:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 484:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 484:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 484:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 484:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 484:18]
  wire  metaArray_clock; // @[Cache.scala 485:25]
  wire  metaArray_reset; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 485:25]
  wire [8:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 485:25]
  wire [16:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 485:25]
  wire [16:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 485:25]
  wire [16:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 485:25]
  wire [16:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 485:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 485:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 485:25]
  wire [8:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 485:25]
  wire [16:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 485:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 485:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 485:25]
  wire  dataArray_clock; // @[Cache.scala 486:25]
  wire  dataArray_reset; // @[Cache.scala 486:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 486:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 486:25]
  wire [11:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 486:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 486:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 486:25]
  wire [11:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 486:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 486:25]
  wire [11:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 486:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 486:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 486:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 495:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 495:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 495:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 495:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 495:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 495:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 495:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 495:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 495:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 495:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 495:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 495:19]
  wire  arb_io_out_ready; // @[Cache.scala 495:19]
  wire  arb_io_out_valid; // @[Cache.scala 495:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 495:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 495:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 495:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 495:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 495:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : REG; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_req_addr; // @[Reg.scala 15:16]
  reg [3:0] r_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_req_wdata; // @[Reg.scala 15:16]
  reg  REG_1; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : REG_1; // @[Pipeline.scala 24:24 25:{25,33}]
  wire  _T_5 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = s2_io_out_valid & s3_io_in_ready | _GEN_8; // @[Pipeline.scala 26:{38,46}]
  reg [31:0] r_1_req_addr; // @[Reg.scala 15:16]
  reg [3:0] r_1_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] r_1_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] r_1_req_wdata; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_0_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_0_dirty; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_1_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_1_dirty; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_2_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_2_dirty; // @[Reg.scala 15:16]
  reg [16:0] r_1_metas_3_tag; // @[Reg.scala 15:16]
  reg  r_1_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] r_1_datas_3_data; // @[Reg.scala 15:16]
  reg  r_1_hit; // @[Reg.scala 15:16]
  reg [3:0] r_1_waymask; // @[Reg.scala 15:16]
  reg  r_1_mmio; // @[Reg.scala 15:16]
  reg  r_1_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] r_1_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] r_1_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_11 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  CacheStage1_2 s1 ( // @[Cache.scala 482:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2_2 s2 ( // @[Cache.scala 483:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3_2 s3 ( // @[Cache.scala 484:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1)
  );
  SRAMTemplateWithArbiter_4 metaArray ( // @[Cache.scala 485:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_5 dataArray ( // @[Cache.scala 486:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 495:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 496:28]
  assign io_in_resp_valid = s3_io_out_valid & _T_11 ? 1'h0 : s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 512:26]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 506:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 506:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 508:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 508:14]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 498:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 498:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 498:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 498:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 498:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 530:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 530:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 531:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 531:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = r_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = r_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = r_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = r_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 537:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 537:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 538:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 538:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 540:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 540:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 539:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 539:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_1; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = r_1_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = r_1_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = r_1_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = r_1_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = r_1_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = r_1_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = r_1_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = r_1_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = r_1_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = r_1_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = r_1_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = r_1_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = r_1_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = r_1_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = r_1_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = r_1_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = r_1_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = r_1_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = r_1_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = r_1_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = r_1_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = r_1_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 532:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 532:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 508:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 508:14]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 530:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 530:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 534:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 534:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 531:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 531:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 532:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 532:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 535:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 535:18]
  assign arb_io_in_0_valid = 1'h0; // @[Cache.scala 520:24]
  assign arb_io_in_0_bits_addr = 32'h0; // @[Cache.scala 517:19 SimpleBus.scala 64:15]
  assign arb_io_in_0_bits_size = 3'h0; // @[Cache.scala 517:19 SimpleBus.scala 66:15]
  assign arb_io_in_0_bits_cmd = 4'h0; // @[Cache.scala 517:19 SimpleBus.scala 65:14]
  assign arb_io_in_0_bits_wmask = 8'h0; // @[Cache.scala 517:19 SimpleBus.scala 68:16]
  assign arb_io_in_0_bits_wdata = 64'h0; // @[Cache.scala 517:19 SimpleBus.scala 67:16]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 496:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 496:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 498:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG <= _GEN_1;
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_cmd <= s1_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wmask <= s1_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      r_req_wdata <= s1_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_1 <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG_1 <= _GEN_9;
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_cmd <= s2_io_out_bits_req_cmd; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wmask <= s2_io_out_bits_req_wmask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_req_wdata <= s2_io_out_bits_req_wdata; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_hit <= s2_io_out_bits_hit; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 16:23]
    end
    if (_T_5) begin // @[Reg.scala 16:19]
      r_1_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_req_cmd = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  r_req_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  r_req_wdata = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_1_req_addr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  r_1_req_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  r_1_req_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  r_1_req_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  r_1_metas_0_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  r_1_metas_0_dirty = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_1_metas_1_tag = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  r_1_metas_1_dirty = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_1_metas_2_tag = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  r_1_metas_2_dirty = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_metas_3_tag = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  r_1_metas_3_dirty = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  r_1_datas_0_data = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  r_1_datas_1_data = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  r_1_datas_2_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  r_1_datas_3_data = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  r_1_hit = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_1_waymask = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  r_1_mmio = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_1_isForwardData = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  r_1_forwardData_data_data = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  r_1_forwardData_waymask = _RAND_27[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusAddressMapper(
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [3:0]  io_out_req_bits_cmd,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
  assign io_in_req_ready = io_out_req_ready; // @[AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = {4'h8,io_in_req_bits_addr[27:0]}; // @[Cat.scala 30:58]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[AddressMapper.scala 31:10]
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  output [2:0]  io_out_awprot,
  output        io_out_awid,
  output        io_out_awuser,
  output [7:0]  io_out_awlen,
  output [2:0]  io_out_awsize,
  output [1:0]  io_out_awburst,
  output        io_out_awlock,
  output [3:0]  io_out_awcache,
  output [3:0]  io_out_awqos,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output        io_out_wlast,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output [2:0]  io_out_arprot,
  output        io_out_arid,
  output        io_out_aruser,
  output [7:0]  io_out_arlen,
  output [2:0]  io_out_arsize,
  output [1:0]  io_out_arburst,
  output        io_out_arlock,
  output [3:0]  io_out_arcache,
  output [3:0]  io_out_arqos,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata,
  input         io_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_rlast ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_17 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_13 & _T_17 & io_out_wlast | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_wlast; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_28 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_36 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_31 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_awprot = io_out_arprot; // @[ToAXI4.scala 182:6]
  assign io_out_awid = io_out_arid; // @[ToAXI4.scala 182:6]
  assign io_out_awuser = io_out_aruser; // @[ToAXI4.scala 182:6]
  assign io_out_awlen = io_out_arlen; // @[ToAXI4.scala 182:6]
  assign io_out_awsize = io_out_arsize; // @[ToAXI4.scala 182:6]
  assign io_out_awburst = io_out_arburst; // @[ToAXI4.scala 182:6]
  assign io_out_awlock = io_out_arlock; // @[ToAXI4.scala 182:6]
  assign io_out_awcache = io_out_arcache; // @[ToAXI4.scala 182:6]
  assign io_out_awqos = io_out_arqos; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_31 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wlast = _T_9 | _T_10; // @[ToAXI4.scala 177:54]
  assign io_out_arvalid = io_in_req_valid & _T_28; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_arprot = 3'h1; // @[ToAXI4.scala 159:12]
  assign io_out_arid = 1'h0; // @[ToAXI4.scala 168:24]
  assign io_out_aruser = 1'h0; // @[ToAXI4.scala 176:24]
  assign io_out_arlen = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:24]
  assign io_out_arsize = 3'h3; // @[ToAXI4.scala 170:24]
  assign io_out_arburst = 2'h2; // @[ToAXI4.scala 171:24]
  assign io_out_arlock = 1'h0; // @[ToAXI4.scala 173:24]
  assign io_out_arcache = 4'h0; // @[ToAXI4.scala 174:24]
  assign io_out_arqos = 4'h0; // @[ToAXI4.scala 175:24]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_23) begin // @[Reg.scala 16:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [2:0]  io_out_0_req_bits_size,
  output [3:0]  io_out_0_req_bits_cmd,
  output [7:0]  io_out_0_req_bits_wmask,
  output [63:0] io_out_0_req_bits_wdata,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [3:0]  io_out_0_resp_bits_cmd,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [3:0]  io_out_1_req_bits_cmd,
  output [7:0]  io_out_1_req_bits_wmask,
  output [63:0] io_out_1_req_bits_wdata,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_out_2_req_ready,
  output        io_out_2_req_valid,
  output [31:0] io_out_2_req_bits_addr,
  output [3:0]  io_out_2_req_bits_cmd,
  output [7:0]  io_out_2_req_bits_wmask,
  output [63:0] io_out_2_req_bits_wdata,
  output        io_out_2_resp_ready,
  input         io_out_2_resp_valid,
  input  [63:0] io_out_2_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[Crossbar.scala 31:22]
  wire  outSelVec_0 = io_in_req_bits_addr >= 32'h40600000 & io_in_req_bits_addr < 32'h41600000; // @[Crossbar.scala 36:34]
  wire  outSelVec_1 = io_in_req_bits_addr >= 32'h38000000 & io_in_req_bits_addr < 32'h38010000; // @[Crossbar.scala 36:34]
  wire  outSelVec_2 = io_in_req_bits_addr >= 32'h3c000000 & io_in_req_bits_addr < 32'h40000000; // @[Crossbar.scala 36:34]
  wire [1:0] _T_9 = outSelVec_1 ? 2'h1 : 2'h2; // @[Mux.scala 47:69]
  wire [1:0] outSelIdx = outSelVec_0 ? 2'h0 : _T_9; // @[Mux.scala 47:69]
  wire  _GEN_1 = 2'h1 == outSelIdx ? io_out_1_req_ready : io_out_0_req_ready; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_2 = 2'h2 == outSelIdx ? io_out_2_req_ready : _GEN_1; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_4 = 2'h1 == outSelIdx ? io_out_1_req_valid : io_out_0_req_valid; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_5 = 2'h2 == outSelIdx ? io_out_2_req_valid : _GEN_4; // @[Decoupled.scala 40:{37,37}]
  wire  _T_10 = _GEN_2 & _GEN_5; // @[Decoupled.scala 40:37]
  wire  _T_11 = state == 2'h0; // @[Crossbar.scala 39:72]
  wire  _T_12 = _T_10 & state == 2'h0; // @[Crossbar.scala 39:62]
  reg [1:0] outSelIdxResp; // @[Reg.scala 15:16]
  wire [2:0] _T_13 = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[Crossbar.scala 41:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_T_13); // @[Crossbar.scala 41:40]
  wire  _T_22 = io_in_req_valid & &_T_13; // @[Crossbar.scala 43:71]
  wire  _GEN_10 = 2'h1 == outSelIdxResp ? io_out_1_resp_ready : io_out_0_resp_ready; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_11 = 2'h2 == outSelIdxResp ? io_out_2_resp_ready : _GEN_10; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_13 = 2'h1 == outSelIdxResp ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Decoupled.scala 40:{37,37}]
  wire  _GEN_14 = 2'h2 == outSelIdxResp ? io_out_2_resp_valid : _GEN_13; // @[Decoupled.scala 40:{37,37}]
  wire  _T_48 = _GEN_11 & _GEN_14; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_16 = io_in_resp_valid ? 2'h0 : state; // @[Crossbar.scala 31:22 64:{43,51}]
  wire [63:0] _GEN_21 = 2'h1 == outSelIdxResp ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Crossbar.scala 68:{19,19}]
  wire [3:0] _GEN_24 = 2'h1 == outSelIdxResp ? 4'h6 : io_out_0_resp_bits_cmd; // @[Crossbar.scala 68:{19,19}]
  assign io_in_req_ready = _GEN_2 | reqInvalidAddr; // @[Crossbar.scala 71:39]
  assign io_in_resp_valid = _T_48 | state == 2'h2; // @[Crossbar.scala 67:46]
  assign io_in_resp_bits_cmd = 2'h2 == outSelIdxResp ? 4'h6 : _GEN_24; // @[Crossbar.scala 68:{19,19}]
  assign io_in_resp_bits_rdata = 2'h2 == outSelIdxResp ? io_out_2_resp_bits_rdata : _GEN_21; // @[Crossbar.scala 68:{19,19}]
  assign io_out_0_req_valid = outSelVec_0 & (io_in_req_valid & _T_11); // @[Crossbar.scala 54:22]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_0_resp_ready = 2'h0 == outSelIdxResp | outSelVec_0; // @[Crossbar.scala 55:18 70:{25,25}]
  assign io_out_1_req_valid = outSelVec_1 & (io_in_req_valid & _T_11); // @[Crossbar.scala 54:22]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_1_resp_ready = 2'h1 == outSelIdxResp | outSelVec_1; // @[Crossbar.scala 55:18 70:{25,25}]
  assign io_out_2_req_valid = outSelVec_2 & (io_in_req_valid & _T_11); // @[Crossbar.scala 54:22]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_2_resp_ready = 2'h2 == outSelIdxResp | outSelVec_2; // @[Crossbar.scala 55:18 70:{25,25}]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 31:22]
      state <= 2'h0; // @[Crossbar.scala 31:22]
    end else if (2'h0 == state) begin // @[Crossbar.scala 58:18]
      if (reqInvalidAddr) begin // @[Crossbar.scala 61:29]
        state <= 2'h2; // @[Crossbar.scala 61:37]
      end else if (_T_10) begin // @[Crossbar.scala 60:32]
        state <= 2'h1; // @[Crossbar.scala 60:40]
      end
    end else if (2'h1 == state) begin // @[Crossbar.scala 58:18]
      if (_T_48) begin // @[Crossbar.scala 63:49]
        state <= 2'h0; // @[Crossbar.scala 63:57]
      end
    end else if (2'h2 == state) begin // @[Crossbar.scala 58:18]
      state <= _GEN_16;
    end
    if (_T_12) begin // @[Reg.scala 16:19]
      if (outSelVec_0) begin // @[Mux.scala 47:69]
        outSelIdxResp <= 2'h0;
      end else if (outSelVec_1) begin // @[Mux.scala 47:69]
        outSelIdxResp <= 2'h1;
      end else begin
        outSelIdxResp <= 2'h2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_22 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!(io.in.req.valid && outSelVec.asUInt.andR), \"address decode error, bad addr = 0x%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_22 | reset)) begin
          $fatal; // @[Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelIdxResp = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  output [2:0]  io_out_awprot,
  output        io_out_awid,
  output        io_out_awuser,
  output [7:0]  io_out_awlen,
  output [2:0]  io_out_awsize,
  output [1:0]  io_out_awburst,
  output        io_out_awlock,
  output [3:0]  io_out_awcache,
  output [3:0]  io_out_awqos,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_wlast,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output [2:0]  io_out_arprot,
  output        io_out_arid,
  output        io_out_aruser,
  output [7:0]  io_out_arlen,
  output [2:0]  io_out_arsize,
  output [1:0]  io_out_arburst,
  output        io_out_arlock,
  output [3:0]  io_out_arcache,
  output [3:0]  io_out_arqos,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata,
  input         io_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_rlast ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_17 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_13 & _T_17 & io_out_wlast | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_wlast; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_28 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_36 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_31 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_awprot = io_out_arprot; // @[ToAXI4.scala 182:6]
  assign io_out_awid = io_out_arid; // @[ToAXI4.scala 182:6]
  assign io_out_awuser = io_out_aruser; // @[ToAXI4.scala 182:6]
  assign io_out_awlen = io_out_arlen; // @[ToAXI4.scala 182:6]
  assign io_out_awsize = io_out_arsize; // @[ToAXI4.scala 182:6]
  assign io_out_awburst = io_out_arburst; // @[ToAXI4.scala 182:6]
  assign io_out_awlock = io_out_arlock; // @[ToAXI4.scala 182:6]
  assign io_out_awcache = io_out_arcache; // @[ToAXI4.scala 182:6]
  assign io_out_awqos = io_out_arqos; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_31 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_wlast = _T_9 | _T_10; // @[ToAXI4.scala 177:54]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_28; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_arprot = 3'h1; // @[ToAXI4.scala 159:12]
  assign io_out_arid = 1'h0; // @[ToAXI4.scala 168:24]
  assign io_out_aruser = 1'h0; // @[ToAXI4.scala 176:24]
  assign io_out_arlen = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:24]
  assign io_out_arsize = io_in_req_bits_size; // @[ToAXI4.scala 170:24]
  assign io_out_arburst = 2'h1; // @[ToAXI4.scala 171:24]
  assign io_out_arlock = 1'h0; // @[ToAXI4.scala 173:24]
  assign io_out_arcache = 4'h0; // @[ToAXI4.scala 174:24]
  assign io_out_arqos = 4'h0; // @[ToAXI4.scala 175:24]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_23) begin // @[Reg.scala 16:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  output        io__extra_mtip,
  output        io__extra_msip,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _T_9 = io__in_wstrb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_11 = io__in_wstrb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_13 = io__in_wstrb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_15 = io__in_wstrb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_17 = io__in_wstrb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_19 = io__in_wstrb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_21 = io__in_wstrb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_23 = io__in_wstrb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] fullMask = {_T_23,_T_21,_T_19,_T_17,_T_15,_T_13,_T_11,_T_9}; // @[Cat.scala 30:58]
  wire  _T_24 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_25 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_25 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_25 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  reg [63:0] mtime; // @[AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[AXI4CLINT.scala 34:21]
  reg [15:0] freq; // @[AXI4CLINT.scala 37:21]
  reg [15:0] inc; // @[AXI4CLINT.scala 38:20]
  reg [15:0] cnt; // @[AXI4CLINT.scala 40:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[AXI4CLINT.scala 41:21]
  wire  tick = nextCnt == freq; // @[AXI4CLINT.scala 43:23]
  wire [63:0] _GEN_14 = {{48'd0}, inc}; // @[AXI4CLINT.scala 44:32]
  wire [63:0] _T_49 = mtime + _GEN_14; // @[AXI4CLINT.scala 44:32]
  wire  _T_78 = 16'h0 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_79 = 16'h8000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_80 = 16'hbff8 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_81 = 16'h8008 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_82 = 16'h4000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_83 = _T_78 ? msip : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_84 = _T_79 ? freq : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_85 = _T_80 ? mtime : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_86 = _T_81 ? inc : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_87 = _T_82 ? mtimecmp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_15 = {{48'd0}, _T_84}; // @[Mux.scala 27:72]
  wire [63:0] _T_88 = _T_83 | _GEN_15; // @[Mux.scala 27:72]
  wire [63:0] _T_89 = _T_88 | _T_85; // @[Mux.scala 27:72]
  wire [63:0] _GEN_16 = {{48'd0}, _T_86}; // @[Mux.scala 27:72]
  wire [63:0] _T_90 = _T_89 | _GEN_16; // @[Mux.scala 27:72]
  wire [63:0] _T_94 = io__in_wdata & fullMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_95 = ~fullMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_96 = msip & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_97 = _T_94 | _T_96; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_17 = {{48'd0}, freq}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_102 = _GEN_17 & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_103 = _T_94 | _T_102; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_10 = _T_42 & io__in_awaddr[15:0] == 16'h8000 ? _T_103 : {{48'd0}, freq}; // @[RegMap.scala 32:{48,52} AXI4CLINT.scala 37:21]
  wire [63:0] _T_108 = mtime & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_109 = _T_94 | _T_108; // @[BitUtils.scala 32:25]
  wire [63:0] _T_114 = _GEN_14 & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_115 = _T_94 | _T_114; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_12 = _T_42 & io__in_awaddr[15:0] == 16'h8008 ? _T_115 : {{48'd0}, inc}; // @[RegMap.scala 32:{48,52} AXI4CLINT.scala 38:20]
  wire [63:0] _T_120 = mtimecmp & _T_95; // @[BitUtils.scala 32:36]
  wire [63:0] _T_121 = _T_94 | _T_120; // @[BitUtils.scala 32:25]
  reg  REG_3; // @[AXI4CLINT.scala 64:31]
  reg  REG_4; // @[AXI4CLINT.scala 65:31]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io__in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io__in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = _T_90 | _T_87; // @[Mux.scala 27:72]
  assign io__extra_mtip = REG_3; // @[AXI4CLINT.scala 64:21]
  assign io__extra_msip = REG_4; // @[AXI4CLINT.scala 65:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    if (reset) begin // @[AXI4CLINT.scala 32:22]
      mtime <= 64'h0; // @[AXI4CLINT.scala 32:22]
    end else if (_T_42 & io__in_awaddr[15:0] == 16'hbff8) begin // @[RegMap.scala 32:48]
      mtime <= _T_109; // @[RegMap.scala 32:52]
    end else if (tick) begin // @[AXI4CLINT.scala 44:15]
      mtime <= _T_49; // @[AXI4CLINT.scala 44:23]
    end
    if (reset) begin // @[AXI4CLINT.scala 33:25]
      mtimecmp <= 64'h0; // @[AXI4CLINT.scala 33:25]
    end else if (_T_42 & io__in_awaddr[15:0] == 16'h4000) begin // @[RegMap.scala 32:48]
      mtimecmp <= _T_121; // @[RegMap.scala 32:52]
    end
    if (reset) begin // @[AXI4CLINT.scala 34:21]
      msip <= 64'h0; // @[AXI4CLINT.scala 34:21]
    end else if (_T_42 & io__in_awaddr[15:0] == 16'h0) begin // @[RegMap.scala 32:48]
      msip <= _T_97; // @[RegMap.scala 32:52]
    end
    if (reset) begin // @[AXI4CLINT.scala 37:21]
      freq <= 16'h28; // @[AXI4CLINT.scala 37:21]
    end else begin
      freq <= _GEN_10[15:0];
    end
    if (reset) begin // @[AXI4CLINT.scala 38:20]
      inc <= 16'h1; // @[AXI4CLINT.scala 38:20]
    end else begin
      inc <= _GEN_12[15:0];
    end
    if (reset) begin // @[AXI4CLINT.scala 40:20]
      cnt <= 16'h0; // @[AXI4CLINT.scala 40:20]
    end else if (nextCnt < freq) begin // @[AXI4CLINT.scala 42:13]
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    REG_3 <= mtime >= mtimecmp; // @[AXI4CLINT.scala 64:38]
    REG_4 <= msip != 64'h0; // @[AXI4CLINT.scala 65:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  freq = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  inc = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  REG_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_4 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBus2AXI4Converter_2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[ToAXI4.scala 151:20]
  wire  _T_8 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_8 | awAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_12 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_8 & _T_12 | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _GEN_2 = _T_12 | wAck; // @[StopWatch.scala 24:20 30:{20,24}]
  wire  _T_18 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_23 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_26 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_31 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_31 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_26 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_26 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_23; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_18) begin // @[Reg.scala 16:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 16:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(toAXI4Lite | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(toAXI4Lite | reset)) begin
          $fatal; // @[ToAXI4.scala 153:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  input  [2:0]  io__extra_intrVec,
  output        io__extra_meip_0,
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _T_24 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_25 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_25 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_25 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  reg [31:0] priority_0; // @[AXI4PLIC.scala 37:39]
  reg [31:0] priority_1; // @[AXI4PLIC.scala 37:39]
  reg [31:0] priority_2; // @[AXI4PLIC.scala 37:39]
  reg  pending_0_1; // @[AXI4PLIC.scala 43:46]
  reg  pending_0_2; // @[AXI4PLIC.scala 43:46]
  reg  pending_0_3; // @[AXI4PLIC.scala 43:46]
  wire [31:0] _T_45 = {16'h0,8'h0,4'h0,pending_0_3,pending_0_2,pending_0_1,1'h0}; // @[Cat.scala 30:58]
  reg [31:0] enable_0_0; // @[AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[AXI4PLIC.scala 53:40]
  reg  inHandle_1; // @[AXI4PLIC.scala 58:25]
  reg  inHandle_2; // @[AXI4PLIC.scala 58:25]
  reg  inHandle_3; // @[AXI4PLIC.scala 58:25]
  reg [31:0] claimCompletion_0; // @[AXI4PLIC.scala 64:46]
  wire  _GEN_13 = _T_25 & io__in_araddr[25:0] == 26'h200004 ? 2'h1 == claimCompletion_0[1:0] | inHandle_1 :
    inHandle_1; // @[AXI4PLIC.scala 58:25 68:59]
  wire  _GEN_14 = _T_25 & io__in_araddr[25:0] == 26'h200004 ? 2'h2 == claimCompletion_0[1:0] | inHandle_2 :
    inHandle_2; // @[AXI4PLIC.scala 58:25 68:59]
  wire  _GEN_15 = _T_25 & io__in_araddr[25:0] == 26'h200004 ? 2'h3 == claimCompletion_0[1:0] | inHandle_3 :
    inHandle_3; // @[AXI4PLIC.scala 58:25 68:59]
  wire  _GEN_16 = io__extra_intrVec[0] | pending_0_1; // @[AXI4PLIC.scala 75:{17,45} 43:46]
  wire  _GEN_18 = io__extra_intrVec[1] | pending_0_2; // @[AXI4PLIC.scala 75:{17,45} 43:46]
  wire  _GEN_20 = io__extra_intrVec[2] | pending_0_3; // @[AXI4PLIC.scala 75:{17,45} 43:46]
  wire [31:0] _T_54 = _T_45 & enable_0_0; // @[AXI4PLIC.scala 81:31]
  wire [4:0] _T_88 = _T_54[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:69]
  wire [4:0] _T_89 = _T_54[29] ? 5'h1d : _T_88; // @[Mux.scala 47:69]
  wire [4:0] _T_90 = _T_54[28] ? 5'h1c : _T_89; // @[Mux.scala 47:69]
  wire [4:0] _T_91 = _T_54[27] ? 5'h1b : _T_90; // @[Mux.scala 47:69]
  wire [4:0] _T_92 = _T_54[26] ? 5'h1a : _T_91; // @[Mux.scala 47:69]
  wire [4:0] _T_93 = _T_54[25] ? 5'h19 : _T_92; // @[Mux.scala 47:69]
  wire [4:0] _T_94 = _T_54[24] ? 5'h18 : _T_93; // @[Mux.scala 47:69]
  wire [4:0] _T_95 = _T_54[23] ? 5'h17 : _T_94; // @[Mux.scala 47:69]
  wire [4:0] _T_96 = _T_54[22] ? 5'h16 : _T_95; // @[Mux.scala 47:69]
  wire [4:0] _T_97 = _T_54[21] ? 5'h15 : _T_96; // @[Mux.scala 47:69]
  wire [4:0] _T_98 = _T_54[20] ? 5'h14 : _T_97; // @[Mux.scala 47:69]
  wire [4:0] _T_99 = _T_54[19] ? 5'h13 : _T_98; // @[Mux.scala 47:69]
  wire [4:0] _T_100 = _T_54[18] ? 5'h12 : _T_99; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = _T_54[17] ? 5'h11 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = _T_54[16] ? 5'h10 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = _T_54[15] ? 5'hf : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = _T_54[14] ? 5'he : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = _T_54[13] ? 5'hd : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = _T_54[12] ? 5'hc : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = _T_54[11] ? 5'hb : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = _T_54[10] ? 5'ha : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = _T_54[9] ? 5'h9 : _T_108; // @[Mux.scala 47:69]
  wire [4:0] _T_110 = _T_54[8] ? 5'h8 : _T_109; // @[Mux.scala 47:69]
  wire [4:0] _T_111 = _T_54[7] ? 5'h7 : _T_110; // @[Mux.scala 47:69]
  wire [4:0] _T_112 = _T_54[6] ? 5'h6 : _T_111; // @[Mux.scala 47:69]
  wire [4:0] _T_113 = _T_54[5] ? 5'h5 : _T_112; // @[Mux.scala 47:69]
  wire [4:0] _T_114 = _T_54[4] ? 5'h4 : _T_113; // @[Mux.scala 47:69]
  wire [4:0] _T_115 = _T_54[3] ? 5'h3 : _T_114; // @[Mux.scala 47:69]
  wire [4:0] _T_116 = _T_54[2] ? 5'h2 : _T_115; // @[Mux.scala 47:69]
  wire [4:0] _T_117 = _T_54[1] ? 5'h1 : _T_116; // @[Mux.scala 47:69]
  wire [4:0] _T_118 = _T_54[0] ? 5'h0 : _T_117; // @[Mux.scala 47:69]
  wire [4:0] _T_119 = _T_54 == 32'h0 ? 5'h0 : _T_118; // @[AXI4PLIC.scala 82:13]
  wire [7:0] _T_124 = io__in_wstrb >> io__in_awaddr[2:0]; // @[AXI4PLIC.scala 89:78]
  wire [7:0] _T_134 = _T_124[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_136 = _T_124[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_138 = _T_124[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_140 = _T_124[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_142 = _T_124[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_144 = _T_124[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_146 = _T_124[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_148 = _T_124[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_149 = {_T_148,_T_146,_T_144,_T_142,_T_140,_T_138,_T_136,_T_134}; // @[Cat.scala 30:58]
  wire  _T_150 = 26'hc == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_151 = 26'h1000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_152 = 26'h2000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_153 = 26'h8 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_154 = 26'h200004 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_155 = 26'h4 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_156 = 26'h200000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_157 = _T_150 ? priority_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_158 = _T_151 ? _T_45 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_159 = _T_152 ? enable_0_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_160 = _T_153 ? priority_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_161 = _T_154 ? claimCompletion_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_162 = _T_155 ? priority_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_163 = _T_156 ? threshold_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_164 = _T_157 | _T_158; // @[Mux.scala 27:72]
  wire [31:0] _T_165 = _T_164 | _T_159; // @[Mux.scala 27:72]
  wire [31:0] _T_166 = _T_165 | _T_160; // @[Mux.scala 27:72]
  wire [31:0] _T_167 = _T_166 | _T_161; // @[Mux.scala 27:72]
  wire [31:0] _T_168 = _T_167 | _T_162; // @[Mux.scala 27:72]
  wire [31:0] rdata = _T_168 | _T_163; // @[Mux.scala 27:72]
  wire [63:0] _T_172 = io__in_wdata & _T_149; // @[BitUtils.scala 32:13]
  wire [63:0] _T_173 = ~_T_149; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_40 = {{32'd0}, priority_2}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_174 = _GEN_40 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_175 = _T_172 | _T_174; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_22 = _T_42 & io__in_awaddr[25:0] == 26'hc ? _T_175 : {{32'd0}, priority_2}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 37:39]
  wire [63:0] _GEN_41 = {{32'd0}, enable_0_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_180 = _GEN_41 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_181 = _T_172 | _T_180; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_23 = _T_42 & io__in_awaddr[25:0] == 26'h2000 ? _T_181 : {{32'd0}, enable_0_0}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 48:64]
  wire [63:0] _GEN_42 = {{32'd0}, priority_1}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_186 = _GEN_42 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_187 = _T_172 | _T_186; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_24 = _T_42 & io__in_awaddr[25:0] == 26'h8 ? _T_187 : {{32'd0}, priority_1}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 37:39]
  wire [63:0] _GEN_43 = {{32'd0}, claimCompletion_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_192 = _GEN_43 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_193 = _T_172 | _T_192; // @[BitUtils.scala 32:25]
  wire [4:0] _GEN_33 = _T_42 & io__in_awaddr[25:0] == 26'h200004 ? 5'h0 : _T_119; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 82:7]
  wire [63:0] _GEN_44 = {{32'd0}, priority_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_200 = _GEN_44 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_201 = _T_172 | _T_200; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_34 = _T_42 & io__in_awaddr[25:0] == 26'h4 ? _T_201 : {{32'd0}, priority_0}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 37:39]
  wire [63:0] _GEN_45 = {{32'd0}, threshold_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_206 = _GEN_45 & _T_173; // @[BitUtils.scala 32:36]
  wire [63:0] _T_207 = _T_172 | _T_206; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_35 = _T_42 & io__in_awaddr[25:0] == 26'h200000 ? _T_207 : {{32'd0}, threshold_0}; // @[RegMap.scala 32:{48,52} AXI4PLIC.scala 53:40]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io__in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io__in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = {rdata,rdata}; // @[Cat.scala 30:58]
  assign io__extra_meip_0 = claimCompletion_0 != 32'h0; // @[AXI4PLIC.scala 93:87]
  assign io_extra_meip_0 = io__extra_meip_0;
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    priority_0 <= _GEN_34[31:0];
    priority_1 <= _GEN_24[31:0];
    priority_2 <= _GEN_22[31:0];
    if (reset) begin // @[AXI4PLIC.scala 43:46]
      pending_0_1 <= 1'h0; // @[AXI4PLIC.scala 43:46]
    end else if (inHandle_1) begin // @[AXI4PLIC.scala 76:25]
      pending_0_1 <= 1'h0; // @[AXI4PLIC.scala 76:53]
    end else begin
      pending_0_1 <= _GEN_16;
    end
    if (reset) begin // @[AXI4PLIC.scala 43:46]
      pending_0_2 <= 1'h0; // @[AXI4PLIC.scala 43:46]
    end else if (inHandle_2) begin // @[AXI4PLIC.scala 76:25]
      pending_0_2 <= 1'h0; // @[AXI4PLIC.scala 76:53]
    end else begin
      pending_0_2 <= _GEN_18;
    end
    if (reset) begin // @[AXI4PLIC.scala 43:46]
      pending_0_3 <= 1'h0; // @[AXI4PLIC.scala 43:46]
    end else if (inHandle_3) begin // @[AXI4PLIC.scala 76:25]
      pending_0_3 <= 1'h0; // @[AXI4PLIC.scala 76:53]
    end else begin
      pending_0_3 <= _GEN_20;
    end
    if (reset) begin // @[AXI4PLIC.scala 48:64]
      enable_0_0 <= 32'h0; // @[AXI4PLIC.scala 48:64]
    end else begin
      enable_0_0 <= _GEN_23[31:0];
    end
    threshold_0 <= _GEN_35[31:0];
    if (reset) begin // @[AXI4PLIC.scala 58:25]
      inHandle_1 <= 1'h0; // @[AXI4PLIC.scala 58:25]
    end else if (_T_42 & io__in_awaddr[25:0] == 26'h200004) begin // @[RegMap.scala 32:48]
      if (2'h1 == _T_193[1:0]) begin // @[AXI4PLIC.scala 60:27]
        inHandle_1 <= 1'h0; // @[AXI4PLIC.scala 60:27]
      end else begin
        inHandle_1 <= _GEN_13;
      end
    end else begin
      inHandle_1 <= _GEN_13;
    end
    if (reset) begin // @[AXI4PLIC.scala 58:25]
      inHandle_2 <= 1'h0; // @[AXI4PLIC.scala 58:25]
    end else if (_T_42 & io__in_awaddr[25:0] == 26'h200004) begin // @[RegMap.scala 32:48]
      if (2'h2 == _T_193[1:0]) begin // @[AXI4PLIC.scala 60:27]
        inHandle_2 <= 1'h0; // @[AXI4PLIC.scala 60:27]
      end else begin
        inHandle_2 <= _GEN_14;
      end
    end else begin
      inHandle_2 <= _GEN_14;
    end
    if (reset) begin // @[AXI4PLIC.scala 58:25]
      inHandle_3 <= 1'h0; // @[AXI4PLIC.scala 58:25]
    end else if (_T_42 & io__in_awaddr[25:0] == 26'h200004) begin // @[RegMap.scala 32:48]
      if (2'h3 == _T_193[1:0]) begin // @[AXI4PLIC.scala 60:27]
        inHandle_3 <= 1'h0; // @[AXI4PLIC.scala 60:27]
      end else begin
        inHandle_3 <= _GEN_15;
      end
    end else begin
      inHandle_3 <= _GEN_15;
    end
    claimCompletion_0 <= {{27'd0}, _GEN_33};
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  priority_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  priority_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  pending_0_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pending_0_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pending_0_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  enable_0_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  threshold_0 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  inHandle_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inHandle_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inHandle_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  claimCompletion_0 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_awready,
  output        io_mem_awvalid,
  output [31:0] io_mem_awaddr,
  output [2:0]  io_mem_awprot,
  output        io_mem_awid,
  output        io_mem_awuser,
  output [7:0]  io_mem_awlen,
  output [2:0]  io_mem_awsize,
  output [1:0]  io_mem_awburst,
  output        io_mem_awlock,
  output [3:0]  io_mem_awcache,
  output [3:0]  io_mem_awqos,
  input         io_mem_wready,
  output        io_mem_wvalid,
  output [63:0] io_mem_wdata,
  output [7:0]  io_mem_wstrb,
  output        io_mem_wlast,
  output        io_mem_bready,
  input         io_mem_bvalid,
  input  [1:0]  io_mem_bresp,
  input         io_mem_bid,
  input         io_mem_buser,
  input         io_mem_arready,
  output        io_mem_arvalid,
  output [31:0] io_mem_araddr,
  output [2:0]  io_mem_arprot,
  output        io_mem_arid,
  output        io_mem_aruser,
  output [7:0]  io_mem_arlen,
  output [2:0]  io_mem_arsize,
  output [1:0]  io_mem_arburst,
  output        io_mem_arlock,
  output [3:0]  io_mem_arcache,
  output [3:0]  io_mem_arqos,
  output        io_mem_rready,
  input         io_mem_rvalid,
  input  [1:0]  io_mem_rresp,
  input  [63:0] io_mem_rdata,
  input         io_mem_rlast,
  input         io_mem_rid,
  input         io_mem_ruser,
  input         io_mmio_awready,
  output        io_mmio_awvalid,
  output [31:0] io_mmio_awaddr,
  output [2:0]  io_mmio_awprot,
  output        io_mmio_awid,
  output        io_mmio_awuser,
  output [7:0]  io_mmio_awlen,
  output [2:0]  io_mmio_awsize,
  output [1:0]  io_mmio_awburst,
  output        io_mmio_awlock,
  output [3:0]  io_mmio_awcache,
  output [3:0]  io_mmio_awqos,
  input         io_mmio_wready,
  output        io_mmio_wvalid,
  output [63:0] io_mmio_wdata,
  output [7:0]  io_mmio_wstrb,
  output        io_mmio_wlast,
  output        io_mmio_bready,
  input         io_mmio_bvalid,
  input  [1:0]  io_mmio_bresp,
  input         io_mmio_bid,
  input         io_mmio_buser,
  input         io_mmio_arready,
  output        io_mmio_arvalid,
  output [31:0] io_mmio_araddr,
  output [2:0]  io_mmio_arprot,
  output        io_mmio_arid,
  output        io_mmio_aruser,
  output [7:0]  io_mmio_arlen,
  output [2:0]  io_mmio_arsize,
  output [1:0]  io_mmio_arburst,
  output        io_mmio_arlock,
  output [3:0]  io_mmio_arcache,
  output [3:0]  io_mmio_arqos,
  output        io_mmio_rready,
  input         io_mmio_rvalid,
  input  [1:0]  io_mmio_rresp,
  input  [63:0] io_mmio_rdata,
  input         io_mmio_rlast,
  input         io_mmio_rid,
  input         io_mmio_ruser,
  output        io_frontend_awready,
  input         io_frontend_awvalid,
  input  [31:0] io_frontend_awaddr,
  input  [2:0]  io_frontend_awprot,
  input         io_frontend_awid,
  input         io_frontend_awuser,
  input  [7:0]  io_frontend_awlen,
  input  [2:0]  io_frontend_awsize,
  input  [1:0]  io_frontend_awburst,
  input         io_frontend_awlock,
  input  [3:0]  io_frontend_awcache,
  input  [3:0]  io_frontend_awqos,
  output        io_frontend_wready,
  input         io_frontend_wvalid,
  input  [63:0] io_frontend_wdata,
  input  [7:0]  io_frontend_wstrb,
  input         io_frontend_wlast,
  input         io_frontend_bready,
  output        io_frontend_bvalid,
  output [1:0]  io_frontend_bresp,
  output        io_frontend_bid,
  output        io_frontend_buser,
  output        io_frontend_arready,
  input         io_frontend_arvalid,
  input  [31:0] io_frontend_araddr,
  input  [2:0]  io_frontend_arprot,
  input         io_frontend_arid,
  input         io_frontend_aruser,
  input  [7:0]  io_frontend_arlen,
  input  [2:0]  io_frontend_arsize,
  input  [1:0]  io_frontend_arburst,
  input         io_frontend_arlock,
  input  [3:0]  io_frontend_arcache,
  input  [3:0]  io_frontend_arqos,
  input         io_frontend_rready,
  output        io_frontend_rvalid,
  output [1:0]  io_frontend_rresp,
  output [63:0] io_frontend_rdata,
  output        io_frontend_rlast,
  output        io_frontend_rid,
  output        io_frontend_ruser,
  input  [2:0]  io_meip,
  output [38:0] io_ila_WBUpc,
  output        io_ila_WBUvalid,
  output        io_ila_WBUrfWen,
  output [4:0]  io_ila_WBUrfDest,
  output [63:0] io_ila_WBUrfData,
  output [63:0] io_ila_InstrCnt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  nutcore_clock; // @[NutShell.scala 53:23]
  wire  nutcore_reset; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_coh_req_bits_addr; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_mmio_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_frontend_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_frontend_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_frontend_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_perfCnts_2; // @[NutShell.scala 53:23]
  wire [38:0] nutcore_io_in_bits_decode_cf_pc; // @[NutShell.scala 53:23]
  wire [4:0] nutcore_io_wb_rfDest; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[NutShell.scala 53:23]
  wire  nutcore_io_wb_rfWen; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_wb_rfData; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[NutShell.scala 53:23]
  wire  nutcore_io_in_valid_0; // @[NutShell.scala 53:23]
  wire  cohMg_clock; // @[NutShell.scala 54:21]
  wire  cohMg_reset; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_coh_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  xbar_clock; // @[NutShell.scala 55:20]
  wire  xbar_reset; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_0_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  axi2sb_clock; // @[NutShell.scala 61:22]
  wire  axi2sb_reset; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_awready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_awvalid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_awaddr; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_awid; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_awlen; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_awsize; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wvalid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_wdata; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_wstrb; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wlast; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_bready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_bvalid; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_arready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_arvalid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_araddr; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_arid; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_arlen; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_arsize; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rvalid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_rdata; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rlast; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_rid; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_valid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_out_req_bits_addr; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_out_req_bits_size; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_valid; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_resp_bits_cmd; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_resp_bits_rdata; // @[NutShell.scala 61:22]
  wire  Prefetcher_clock; // @[NutShell.scala 73:30]
  wire  Prefetcher_reset; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_in_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_in_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_in_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_in_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_in_bits_wdata; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_out_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_out_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_out_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_out_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_out_bits_wdata; // @[NutShell.scala 73:30]
  wire  Cache_clock; // @[Cache.scala 670:35]
  wire  Cache_reset; // @[Cache.scala 670:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 670:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 670:35]
  wire [2:0] Cache_io_in_req_bits_size; // @[Cache.scala 670:35]
  wire [3:0] Cache_io_in_req_bits_cmd; // @[Cache.scala 670:35]
  wire [7:0] Cache_io_in_req_bits_wmask; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_in_req_bits_wdata; // @[Cache.scala 670:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 670:35]
  wire [3:0] Cache_io_in_resp_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 670:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 670:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 670:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 670:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 670:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 670:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 670:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 670:35]
  wire  memAddrMap_io_in_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  SimpleBus2AXI4Converter_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_awprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awuser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_awlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_awsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_awburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_awcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_awqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wlast; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_arprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_aruser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_arlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_arsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_arburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_arcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_arqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rlast; // @[ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_in_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_0_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  SimpleBus2AXI4Converter_1_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_in_req_bits_size; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_awprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awuser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_awlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_awsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_1_io_out_awburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_awcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_awqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wlast; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_arprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_aruser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_arlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_arsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_1_io_out_arburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_arcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_arqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rlast; // @[ToAXI4.scala 204:24]
  wire  clint_clock; // @[NutShell.scala 113:21]
  wire  clint_reset; // @[NutShell.scala 113:21]
  wire  clint_io__in_awready; // @[NutShell.scala 113:21]
  wire  clint_io__in_awvalid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_awaddr; // @[NutShell.scala 113:21]
  wire  clint_io__in_wready; // @[NutShell.scala 113:21]
  wire  clint_io__in_wvalid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_wdata; // @[NutShell.scala 113:21]
  wire [7:0] clint_io__in_wstrb; // @[NutShell.scala 113:21]
  wire  clint_io__in_bready; // @[NutShell.scala 113:21]
  wire  clint_io__in_bvalid; // @[NutShell.scala 113:21]
  wire  clint_io__in_arready; // @[NutShell.scala 113:21]
  wire  clint_io__in_arvalid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_araddr; // @[NutShell.scala 113:21]
  wire  clint_io__in_rready; // @[NutShell.scala 113:21]
  wire  clint_io__in_rvalid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_rdata; // @[NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[NutShell.scala 113:21]
  wire  SimpleBus2AXI4Converter_2_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_2_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  plic_clock; // @[NutShell.scala 120:20]
  wire  plic_reset; // @[NutShell.scala 120:20]
  wire  plic_io__in_awready; // @[NutShell.scala 120:20]
  wire  plic_io__in_awvalid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_awaddr; // @[NutShell.scala 120:20]
  wire  plic_io__in_wready; // @[NutShell.scala 120:20]
  wire  plic_io__in_wvalid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_wdata; // @[NutShell.scala 120:20]
  wire [7:0] plic_io__in_wstrb; // @[NutShell.scala 120:20]
  wire  plic_io__in_bready; // @[NutShell.scala 120:20]
  wire  plic_io__in_bvalid; // @[NutShell.scala 120:20]
  wire  plic_io__in_arready; // @[NutShell.scala 120:20]
  wire  plic_io__in_arvalid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_araddr; // @[NutShell.scala 120:20]
  wire  plic_io__in_rready; // @[NutShell.scala 120:20]
  wire  plic_io__in_rvalid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_rdata; // @[NutShell.scala 120:20]
  wire [2:0] plic_io__extra_intrVec; // @[NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[NutShell.scala 120:20]
  wire  SimpleBus2AXI4Converter_3_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_3_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_rdata; // @[ToAXI4.scala 204:24]
  reg [2:0] REG; // @[NutShell.scala 122:47]
  reg [2:0] REG_1; // @[NutShell.scala 122:39]
  wire  ilaWBUvalid = nutcore_io_in_valid_0;
  wire  ilaWBUrfWen = nutcore_io_wb_rfWen;
  wire [4:0] ilaWBUrfDest = nutcore_io_wb_rfDest;
  wire [38:0] ilaWBUpc = nutcore_io_in_bits_decode_cf_pc;
  wire [63:0] _WIRE_6 = {{25'd0}, ilaWBUpc};
  wire [63:0] _WIRE_7 = {{63'd0}, ilaWBUvalid};
  wire [63:0] _WIRE_8 = {{63'd0}, ilaWBUrfWen};
  wire [63:0] _WIRE_9 = {{59'd0}, ilaWBUrfDest};
  NutCore nutcore ( // @[NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_req_bits_cmd(nutcore_io_imem_mem_req_bits_cmd),
    .io_imem_mem_req_bits_wdata(nutcore_io_imem_mem_req_bits_wdata),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_cmd(nutcore_io_imem_mem_resp_bits_cmd),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_dmem_coh_req_ready(nutcore_io_dmem_coh_req_ready),
    .io_dmem_coh_req_valid(nutcore_io_dmem_coh_req_valid),
    .io_dmem_coh_req_bits_addr(nutcore_io_dmem_coh_req_bits_addr),
    .io_dmem_coh_req_bits_wdata(nutcore_io_dmem_coh_req_bits_wdata),
    .io_dmem_coh_resp_valid(nutcore_io_dmem_coh_resp_valid),
    .io_dmem_coh_resp_bits_cmd(nutcore_io_dmem_coh_resp_bits_cmd),
    .io_dmem_coh_resp_bits_rdata(nutcore_io_dmem_coh_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(nutcore_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_frontend_req_ready(nutcore_io_frontend_req_ready),
    .io_frontend_req_valid(nutcore_io_frontend_req_valid),
    .io_frontend_req_bits_addr(nutcore_io_frontend_req_bits_addr),
    .io_frontend_req_bits_size(nutcore_io_frontend_req_bits_size),
    .io_frontend_req_bits_cmd(nutcore_io_frontend_req_bits_cmd),
    .io_frontend_req_bits_wmask(nutcore_io_frontend_req_bits_wmask),
    .io_frontend_req_bits_wdata(nutcore_io_frontend_req_bits_wdata),
    .io_frontend_resp_ready(nutcore_io_frontend_resp_ready),
    .io_frontend_resp_valid(nutcore_io_frontend_resp_valid),
    .io_frontend_resp_bits_cmd(nutcore_io_frontend_resp_bits_cmd),
    .io_frontend_resp_bits_rdata(nutcore_io_frontend_resp_bits_rdata),
    .perfCnts_2(nutcore_perfCnts_2),
    .io_in_bits_decode_cf_pc(nutcore_io_in_bits_decode_cf_pc),
    .io_wb_rfDest(nutcore_io_wb_rfDest),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    .io_wb_rfWen(nutcore_io_wb_rfWen),
    .io_wb_rfData(nutcore_io_wb_rfData),
    .io_extra_msip(nutcore_io_extra_msip),
    .io_in_valid_0(nutcore_io_in_valid_0)
  );
  CoherenceManager cohMg ( // @[NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_req_bits_cmd(cohMg_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(cohMg_io_in_req_bits_wdata),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(cohMg_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(cohMg_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(cohMg_io_out_coh_req_ready),
    .io_out_coh_req_valid(cohMg_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(cohMg_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(cohMg_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_ready(cohMg_io_out_coh_resp_ready),
    .io_out_coh_resp_valid(cohMg_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(cohMg_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(cohMg_io_out_coh_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1 xbar ( // @[NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(xbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(xbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(xbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  AXI42SimpleBusConverter axi2sb ( // @[NutShell.scala 61:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset),
    .io_in_awready(axi2sb_io_in_awready),
    .io_in_awvalid(axi2sb_io_in_awvalid),
    .io_in_awaddr(axi2sb_io_in_awaddr),
    .io_in_awid(axi2sb_io_in_awid),
    .io_in_awlen(axi2sb_io_in_awlen),
    .io_in_awsize(axi2sb_io_in_awsize),
    .io_in_wready(axi2sb_io_in_wready),
    .io_in_wvalid(axi2sb_io_in_wvalid),
    .io_in_wdata(axi2sb_io_in_wdata),
    .io_in_wstrb(axi2sb_io_in_wstrb),
    .io_in_wlast(axi2sb_io_in_wlast),
    .io_in_bready(axi2sb_io_in_bready),
    .io_in_bvalid(axi2sb_io_in_bvalid),
    .io_in_arready(axi2sb_io_in_arready),
    .io_in_arvalid(axi2sb_io_in_arvalid),
    .io_in_araddr(axi2sb_io_in_araddr),
    .io_in_arid(axi2sb_io_in_arid),
    .io_in_arlen(axi2sb_io_in_arlen),
    .io_in_arsize(axi2sb_io_in_arsize),
    .io_in_rready(axi2sb_io_in_rready),
    .io_in_rvalid(axi2sb_io_in_rvalid),
    .io_in_rdata(axi2sb_io_in_rdata),
    .io_in_rlast(axi2sb_io_in_rlast),
    .io_in_rid(axi2sb_io_in_rid),
    .io_out_req_ready(axi2sb_io_out_req_ready),
    .io_out_req_valid(axi2sb_io_out_req_valid),
    .io_out_req_bits_addr(axi2sb_io_out_req_bits_addr),
    .io_out_req_bits_size(axi2sb_io_out_req_bits_size),
    .io_out_req_bits_cmd(axi2sb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(axi2sb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(axi2sb_io_out_req_bits_wdata),
    .io_out_resp_ready(axi2sb_io_out_resp_ready),
    .io_out_resp_valid(axi2sb_io_out_resp_valid),
    .io_out_resp_bits_cmd(axi2sb_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(axi2sb_io_out_resp_bits_rdata)
  );
  Prefetcher Prefetcher ( // @[NutShell.scala 73:30]
    .clock(Prefetcher_clock),
    .reset(Prefetcher_reset),
    .io_in_ready(Prefetcher_io_in_ready),
    .io_in_valid(Prefetcher_io_in_valid),
    .io_in_bits_addr(Prefetcher_io_in_bits_addr),
    .io_in_bits_size(Prefetcher_io_in_bits_size),
    .io_in_bits_cmd(Prefetcher_io_in_bits_cmd),
    .io_in_bits_wmask(Prefetcher_io_in_bits_wmask),
    .io_in_bits_wdata(Prefetcher_io_in_bits_wdata),
    .io_out_ready(Prefetcher_io_out_ready),
    .io_out_valid(Prefetcher_io_out_valid),
    .io_out_bits_addr(Prefetcher_io_out_bits_addr),
    .io_out_bits_size(Prefetcher_io_out_bits_size),
    .io_out_bits_cmd(Prefetcher_io_out_bits_cmd),
    .io_out_bits_wmask(Prefetcher_io_out_bits_wmask),
    .io_out_bits_wdata(Prefetcher_io_out_bits_wdata)
  );
  Cache_2 Cache ( // @[Cache.scala 670:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_io_in_req_bits_wdata),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata)
  );
  SimpleBusAddressMapper memAddrMap ( // @[NutShell.scala 93:26]
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter SimpleBus2AXI4Converter ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_clock),
    .reset(SimpleBus2AXI4Converter_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_io_in_req_bits_wdata),
    .io_in_resp_valid(SimpleBus2AXI4Converter_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_io_out_awaddr),
    .io_out_awprot(SimpleBus2AXI4Converter_io_out_awprot),
    .io_out_awid(SimpleBus2AXI4Converter_io_out_awid),
    .io_out_awuser(SimpleBus2AXI4Converter_io_out_awuser),
    .io_out_awlen(SimpleBus2AXI4Converter_io_out_awlen),
    .io_out_awsize(SimpleBus2AXI4Converter_io_out_awsize),
    .io_out_awburst(SimpleBus2AXI4Converter_io_out_awburst),
    .io_out_awlock(SimpleBus2AXI4Converter_io_out_awlock),
    .io_out_awcache(SimpleBus2AXI4Converter_io_out_awcache),
    .io_out_awqos(SimpleBus2AXI4Converter_io_out_awqos),
    .io_out_wready(SimpleBus2AXI4Converter_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_io_out_wdata),
    .io_out_wlast(SimpleBus2AXI4Converter_io_out_wlast),
    .io_out_bvalid(SimpleBus2AXI4Converter_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_io_out_araddr),
    .io_out_arprot(SimpleBus2AXI4Converter_io_out_arprot),
    .io_out_arid(SimpleBus2AXI4Converter_io_out_arid),
    .io_out_aruser(SimpleBus2AXI4Converter_io_out_aruser),
    .io_out_arlen(SimpleBus2AXI4Converter_io_out_arlen),
    .io_out_arsize(SimpleBus2AXI4Converter_io_out_arsize),
    .io_out_arburst(SimpleBus2AXI4Converter_io_out_arburst),
    .io_out_arlock(SimpleBus2AXI4Converter_io_out_arlock),
    .io_out_arcache(SimpleBus2AXI4Converter_io_out_arcache),
    .io_out_arqos(SimpleBus2AXI4Converter_io_out_arqos),
    .io_out_rvalid(SimpleBus2AXI4Converter_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_io_out_rdata),
    .io_out_rlast(SimpleBus2AXI4Converter_io_out_rlast)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_size(mmioXbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_size(mmioXbar_io_out_0_req_bits_size),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_cmd(mmioXbar_io_out_0_resp_bits_cmd),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_1 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_1_clock),
    .reset(SimpleBus2AXI4Converter_1_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_1_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_1_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_1_io_in_req_bits_addr),
    .io_in_req_bits_size(SimpleBus2AXI4Converter_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_1_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_1_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_1_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_1_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_1_io_out_awaddr),
    .io_out_awprot(SimpleBus2AXI4Converter_1_io_out_awprot),
    .io_out_awid(SimpleBus2AXI4Converter_1_io_out_awid),
    .io_out_awuser(SimpleBus2AXI4Converter_1_io_out_awuser),
    .io_out_awlen(SimpleBus2AXI4Converter_1_io_out_awlen),
    .io_out_awsize(SimpleBus2AXI4Converter_1_io_out_awsize),
    .io_out_awburst(SimpleBus2AXI4Converter_1_io_out_awburst),
    .io_out_awlock(SimpleBus2AXI4Converter_1_io_out_awlock),
    .io_out_awcache(SimpleBus2AXI4Converter_1_io_out_awcache),
    .io_out_awqos(SimpleBus2AXI4Converter_1_io_out_awqos),
    .io_out_wready(SimpleBus2AXI4Converter_1_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_1_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_1_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_1_io_out_wstrb),
    .io_out_wlast(SimpleBus2AXI4Converter_1_io_out_wlast),
    .io_out_bready(SimpleBus2AXI4Converter_1_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_1_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_1_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_1_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_1_io_out_araddr),
    .io_out_arprot(SimpleBus2AXI4Converter_1_io_out_arprot),
    .io_out_arid(SimpleBus2AXI4Converter_1_io_out_arid),
    .io_out_aruser(SimpleBus2AXI4Converter_1_io_out_aruser),
    .io_out_arlen(SimpleBus2AXI4Converter_1_io_out_arlen),
    .io_out_arsize(SimpleBus2AXI4Converter_1_io_out_arsize),
    .io_out_arburst(SimpleBus2AXI4Converter_1_io_out_arburst),
    .io_out_arlock(SimpleBus2AXI4Converter_1_io_out_arlock),
    .io_out_arcache(SimpleBus2AXI4Converter_1_io_out_arcache),
    .io_out_arqos(SimpleBus2AXI4Converter_1_io_out_arqos),
    .io_out_rready(SimpleBus2AXI4Converter_1_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_1_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_1_io_out_rdata),
    .io_out_rlast(SimpleBus2AXI4Converter_1_io_out_rlast)
  );
  AXI4CLINT clint ( // @[NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_awready(clint_io__in_awready),
    .io__in_awvalid(clint_io__in_awvalid),
    .io__in_awaddr(clint_io__in_awaddr),
    .io__in_wready(clint_io__in_wready),
    .io__in_wvalid(clint_io__in_wvalid),
    .io__in_wdata(clint_io__in_wdata),
    .io__in_wstrb(clint_io__in_wstrb),
    .io__in_bready(clint_io__in_bready),
    .io__in_bvalid(clint_io__in_bvalid),
    .io__in_arready(clint_io__in_arready),
    .io__in_arvalid(clint_io__in_arvalid),
    .io__in_araddr(clint_io__in_araddr),
    .io__in_rready(clint_io__in_rready),
    .io__in_rvalid(clint_io__in_rvalid),
    .io__in_rdata(clint_io__in_rdata),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_2 SimpleBus2AXI4Converter_2 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_2_clock),
    .reset(SimpleBus2AXI4Converter_2_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_2_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_2_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_2_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_2_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_2_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_2_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_2_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_2_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_2_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_2_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_2_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_2_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_2_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_2_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_2_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_2_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_2_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_2_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_2_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_2_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_2_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_2_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_2_io_out_rdata)
  );
  AXI4PLIC plic ( // @[NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_awready(plic_io__in_awready),
    .io__in_awvalid(plic_io__in_awvalid),
    .io__in_awaddr(plic_io__in_awaddr),
    .io__in_wready(plic_io__in_wready),
    .io__in_wvalid(plic_io__in_wvalid),
    .io__in_wdata(plic_io__in_wdata),
    .io__in_wstrb(plic_io__in_wstrb),
    .io__in_bready(plic_io__in_bready),
    .io__in_bvalid(plic_io__in_bvalid),
    .io__in_arready(plic_io__in_arready),
    .io__in_arvalid(plic_io__in_arvalid),
    .io__in_araddr(plic_io__in_araddr),
    .io__in_rready(plic_io__in_rready),
    .io__in_rvalid(plic_io__in_rvalid),
    .io__in_rdata(plic_io__in_rdata),
    .io__extra_intrVec(plic_io__extra_intrVec),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_2 SimpleBus2AXI4Converter_3 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_3_clock),
    .reset(SimpleBus2AXI4Converter_3_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_3_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_3_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_3_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_3_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_3_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_3_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_3_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_3_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_3_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_3_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_3_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_3_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_3_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_3_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_3_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_3_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_3_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_3_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_3_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_3_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_3_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_3_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_3_io_out_rdata)
  );
  assign io_mem_awvalid = SimpleBus2AXI4Converter_io_out_awvalid; // @[NutShell.scala 95:10]
  assign io_mem_awaddr = SimpleBus2AXI4Converter_io_out_awaddr; // @[NutShell.scala 95:10]
  assign io_mem_awprot = SimpleBus2AXI4Converter_io_out_awprot; // @[NutShell.scala 95:10]
  assign io_mem_awid = SimpleBus2AXI4Converter_io_out_awid; // @[NutShell.scala 95:10]
  assign io_mem_awuser = SimpleBus2AXI4Converter_io_out_awuser; // @[NutShell.scala 95:10]
  assign io_mem_awlen = SimpleBus2AXI4Converter_io_out_awlen; // @[NutShell.scala 95:10]
  assign io_mem_awsize = SimpleBus2AXI4Converter_io_out_awsize; // @[NutShell.scala 95:10]
  assign io_mem_awburst = SimpleBus2AXI4Converter_io_out_awburst; // @[NutShell.scala 95:10]
  assign io_mem_awlock = SimpleBus2AXI4Converter_io_out_awlock; // @[NutShell.scala 95:10]
  assign io_mem_awcache = SimpleBus2AXI4Converter_io_out_awcache; // @[NutShell.scala 95:10]
  assign io_mem_awqos = SimpleBus2AXI4Converter_io_out_awqos; // @[NutShell.scala 95:10]
  assign io_mem_wvalid = SimpleBus2AXI4Converter_io_out_wvalid; // @[NutShell.scala 95:10]
  assign io_mem_wdata = SimpleBus2AXI4Converter_io_out_wdata; // @[NutShell.scala 95:10]
  assign io_mem_wstrb = 8'hff; // @[NutShell.scala 95:10]
  assign io_mem_wlast = SimpleBus2AXI4Converter_io_out_wlast; // @[NutShell.scala 95:10]
  assign io_mem_bready = 1'h1; // @[NutShell.scala 95:10]
  assign io_mem_arvalid = SimpleBus2AXI4Converter_io_out_arvalid; // @[NutShell.scala 95:10]
  assign io_mem_araddr = SimpleBus2AXI4Converter_io_out_araddr; // @[NutShell.scala 95:10]
  assign io_mem_arprot = 3'h1; // @[NutShell.scala 95:10]
  assign io_mem_arid = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_aruser = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_arlen = SimpleBus2AXI4Converter_io_out_arlen; // @[NutShell.scala 95:10]
  assign io_mem_arsize = 3'h3; // @[NutShell.scala 95:10]
  assign io_mem_arburst = 2'h2; // @[NutShell.scala 95:10]
  assign io_mem_arlock = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_arcache = 4'h0; // @[NutShell.scala 95:10]
  assign io_mem_arqos = 4'h0; // @[NutShell.scala 95:10]
  assign io_mem_rready = 1'h1; // @[NutShell.scala 95:10]
  assign io_mmio_awvalid = SimpleBus2AXI4Converter_1_io_out_awvalid; // @[NutShell.scala 110:33]
  assign io_mmio_awaddr = SimpleBus2AXI4Converter_1_io_out_awaddr; // @[NutShell.scala 110:33]
  assign io_mmio_awprot = SimpleBus2AXI4Converter_1_io_out_awprot; // @[NutShell.scala 110:33]
  assign io_mmio_awid = SimpleBus2AXI4Converter_1_io_out_awid; // @[NutShell.scala 110:33]
  assign io_mmio_awuser = SimpleBus2AXI4Converter_1_io_out_awuser; // @[NutShell.scala 110:33]
  assign io_mmio_awlen = SimpleBus2AXI4Converter_1_io_out_awlen; // @[NutShell.scala 110:33]
  assign io_mmio_awsize = SimpleBus2AXI4Converter_1_io_out_awsize; // @[NutShell.scala 110:33]
  assign io_mmio_awburst = SimpleBus2AXI4Converter_1_io_out_awburst; // @[NutShell.scala 110:33]
  assign io_mmio_awlock = SimpleBus2AXI4Converter_1_io_out_awlock; // @[NutShell.scala 110:33]
  assign io_mmio_awcache = SimpleBus2AXI4Converter_1_io_out_awcache; // @[NutShell.scala 110:33]
  assign io_mmio_awqos = SimpleBus2AXI4Converter_1_io_out_awqos; // @[NutShell.scala 110:33]
  assign io_mmio_wvalid = SimpleBus2AXI4Converter_1_io_out_wvalid; // @[NutShell.scala 110:33]
  assign io_mmio_wdata = SimpleBus2AXI4Converter_1_io_out_wdata; // @[NutShell.scala 110:33]
  assign io_mmio_wstrb = SimpleBus2AXI4Converter_1_io_out_wstrb; // @[NutShell.scala 110:33]
  assign io_mmio_wlast = SimpleBus2AXI4Converter_1_io_out_wlast; // @[NutShell.scala 110:33]
  assign io_mmio_bready = SimpleBus2AXI4Converter_1_io_out_bready; // @[NutShell.scala 110:33]
  assign io_mmio_arvalid = SimpleBus2AXI4Converter_1_io_out_arvalid; // @[NutShell.scala 110:33]
  assign io_mmio_araddr = SimpleBus2AXI4Converter_1_io_out_araddr; // @[NutShell.scala 110:33]
  assign io_mmio_arprot = 3'h1; // @[NutShell.scala 110:33]
  assign io_mmio_arid = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_aruser = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arlen = SimpleBus2AXI4Converter_1_io_out_arlen; // @[NutShell.scala 110:33]
  assign io_mmio_arsize = SimpleBus2AXI4Converter_1_io_out_arsize; // @[NutShell.scala 110:33]
  assign io_mmio_arburst = 2'h1; // @[NutShell.scala 110:33]
  assign io_mmio_arlock = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arcache = 4'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arqos = 4'h0; // @[NutShell.scala 110:33]
  assign io_mmio_rready = SimpleBus2AXI4Converter_1_io_out_rready; // @[NutShell.scala 110:33]
  assign io_frontend_awready = axi2sb_io_in_awready; // @[NutShell.scala 62:16]
  assign io_frontend_wready = axi2sb_io_in_wready; // @[NutShell.scala 62:16]
  assign io_frontend_bvalid = axi2sb_io_in_bvalid; // @[NutShell.scala 62:16]
  assign io_frontend_bresp = 2'h0; // @[NutShell.scala 62:16]
  assign io_frontend_bid = 1'h0; // @[NutShell.scala 62:16]
  assign io_frontend_buser = 1'h0; // @[NutShell.scala 62:16]
  assign io_frontend_arready = axi2sb_io_in_arready; // @[NutShell.scala 62:16]
  assign io_frontend_rvalid = axi2sb_io_in_rvalid; // @[NutShell.scala 62:16]
  assign io_frontend_rresp = 2'h0; // @[NutShell.scala 62:16]
  assign io_frontend_rdata = axi2sb_io_in_rdata; // @[NutShell.scala 62:16]
  assign io_frontend_rlast = axi2sb_io_in_rlast; // @[NutShell.scala 62:16]
  assign io_frontend_rid = axi2sb_io_in_rid[0]; // @[NutShell.scala 62:16]
  assign io_frontend_ruser = 1'h0; // @[NutShell.scala 62:16]
  assign io_ila_WBUpc = _WIRE_6[38:0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUvalid = _WIRE_7[0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfWen = _WIRE_8[0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfDest = _WIRE_9[4:0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfData = nutcore_io_wb_rfData; // @[NutShell.scala 132:12]
  assign io_ila_InstrCnt = nutcore_perfCnts_2; // @[NutShell.scala 132:12]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_cmd = cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_coh_req_valid = cohMg_io_out_coh_req_valid; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_addr = cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_wdata = cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 57:23]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 107:18]
  assign nutcore_io_frontend_req_valid = axi2sb_io_out_req_valid; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_addr = axi2sb_io_out_req_bits_addr; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_size = axi2sb_io_out_req_bits_size; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_cmd = axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wmask = axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wdata = axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_resp_ready = axi2sb_io_out_resp_ready; // @[NutShell.scala 63:23]
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_cmd = nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_wdata = nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 58:17]
  assign cohMg_io_out_coh_req_ready = nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_valid = nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_cmd = nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_rdata = nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 57:23]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_cmd = cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wmask = 8'hff; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wdata = cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = 3'h3; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = 8'hff; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 59:17]
  assign xbar_io_out_req_ready = Prefetcher_io_in_ready; // @[NutShell.scala 75:24]
  assign xbar_io_out_resp_valid = Cache_io_in_resp_valid; // @[Cache.scala 676:17 NutShell.scala 74:27]
  assign xbar_io_out_resp_bits_cmd = Cache_io_in_resp_bits_cmd; // @[Cache.scala 676:17 NutShell.scala 74:27]
  assign xbar_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[Cache.scala 676:17 NutShell.scala 74:27]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign axi2sb_io_in_awvalid = io_frontend_awvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awaddr = io_frontend_awaddr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awid = {{17'd0}, io_frontend_awid}; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awlen = io_frontend_awlen; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awsize = io_frontend_awsize; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wvalid = io_frontend_wvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wdata = io_frontend_wdata; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wstrb = io_frontend_wstrb; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wlast = io_frontend_wlast; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_bready = io_frontend_bready; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arvalid = io_frontend_arvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_araddr = io_frontend_araddr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arid = {{17'd0}, io_frontend_arid}; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arlen = io_frontend_arlen; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arsize = io_frontend_arsize; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_rready = io_frontend_rready; // @[NutShell.scala 62:16]
  assign axi2sb_io_out_req_ready = nutcore_io_frontend_req_ready; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_valid = nutcore_io_frontend_resp_valid; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_cmd = nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_rdata = nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 63:23]
  assign Prefetcher_clock = clock;
  assign Prefetcher_reset = reset;
  assign Prefetcher_io_in_valid = xbar_io_out_req_valid; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_addr = xbar_io_out_req_bits_addr; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_size = xbar_io_out_req_bits_size; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_cmd = xbar_io_out_req_bits_cmd; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wmask = xbar_io_out_req_bits_wmask; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wdata = xbar_io_out_req_bits_wdata; // @[NutShell.scala 75:24]
  assign Prefetcher_io_out_ready = Cache_io_in_req_ready; // @[Cache.scala 676:17 NutShell.scala 74:27]
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = Prefetcher_io_out_valid; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_addr = Prefetcher_io_out_bits_addr; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_size = Prefetcher_io_out_bits_size; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_cmd = Prefetcher_io_out_bits_cmd; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_wmask = Prefetcher_io_out_bits_wmask; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_in_req_bits_wdata = Prefetcher_io_out_bits_wdata; // @[NutShell.scala 74:27 76:21]
  assign Cache_io_out_mem_req_ready = memAddrMap_io_in_req_ready; // @[NutShell.scala 71:26 94:20]
  assign Cache_io_out_mem_resp_valid = memAddrMap_io_in_resp_valid; // @[NutShell.scala 71:26 94:20]
  assign Cache_io_out_mem_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 71:26 94:20]
  assign Cache_io_out_mem_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 71:26 94:20]
  assign memAddrMap_io_in_req_valid = Cache_io_out_mem_req_valid; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_in_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutShell.scala 71:26 81:16]
  assign memAddrMap_io_out_req_ready = SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_clock = clock;
  assign SimpleBus2AXI4Converter_reset = reset;
  assign SimpleBus2AXI4Converter_io_in_req_valid = memAddrMap_io_out_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_out_awready = io_mem_awready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_wready = io_mem_wready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_bvalid = io_mem_bvalid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_arready = io_mem_arready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rvalid = io_mem_rvalid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rdata = io_mem_rdata; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rlast = io_mem_rlast; // @[NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_size = nutcore_io_mmio_req_bits_size; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_valid = SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_cmd = SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_req_ready = SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_valid = SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_clock = clock;
  assign SimpleBus2AXI4Converter_1_reset = reset;
  assign SimpleBus2AXI4Converter_1_io_in_req_valid = mmioXbar_io_out_0_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_size = mmioXbar_io_out_0_req_bits_size; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_resp_ready = mmioXbar_io_out_0_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_out_awready = io_mmio_awready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_wready = io_mmio_wready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_bvalid = io_mmio_bvalid; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_arready = io_mmio_arready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rvalid = io_mmio_rvalid; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rdata = io_mmio_rdata; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rlast = io_mmio_rlast; // @[NutShell.scala 110:33]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_awvalid = SimpleBus2AXI4Converter_2_io_out_awvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_awaddr = SimpleBus2AXI4Converter_2_io_out_awaddr; // @[NutShell.scala 114:15]
  assign clint_io__in_wvalid = SimpleBus2AXI4Converter_2_io_out_wvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_wdata = SimpleBus2AXI4Converter_2_io_out_wdata; // @[NutShell.scala 114:15]
  assign clint_io__in_wstrb = SimpleBus2AXI4Converter_2_io_out_wstrb; // @[NutShell.scala 114:15]
  assign clint_io__in_bready = SimpleBus2AXI4Converter_2_io_out_bready; // @[NutShell.scala 114:15]
  assign clint_io__in_arvalid = SimpleBus2AXI4Converter_2_io_out_arvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_araddr = SimpleBus2AXI4Converter_2_io_out_araddr; // @[NutShell.scala 114:15]
  assign clint_io__in_rready = SimpleBus2AXI4Converter_2_io_out_rready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_clock = clock;
  assign SimpleBus2AXI4Converter_2_reset = reset;
  assign SimpleBus2AXI4Converter_2_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_out_awready = clint_io__in_awready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_wready = clint_io__in_wready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_bvalid = clint_io__in_bvalid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_arready = clint_io__in_arready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_rvalid = clint_io__in_rvalid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_rdata = clint_io__in_rdata; // @[NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_awvalid = SimpleBus2AXI4Converter_3_io_out_awvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_awaddr = SimpleBus2AXI4Converter_3_io_out_awaddr; // @[NutShell.scala 121:14]
  assign plic_io__in_wvalid = SimpleBus2AXI4Converter_3_io_out_wvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_wdata = SimpleBus2AXI4Converter_3_io_out_wdata; // @[NutShell.scala 121:14]
  assign plic_io__in_wstrb = SimpleBus2AXI4Converter_3_io_out_wstrb; // @[NutShell.scala 121:14]
  assign plic_io__in_bready = SimpleBus2AXI4Converter_3_io_out_bready; // @[NutShell.scala 121:14]
  assign plic_io__in_arvalid = SimpleBus2AXI4Converter_3_io_out_arvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_araddr = SimpleBus2AXI4Converter_3_io_out_araddr; // @[NutShell.scala 121:14]
  assign plic_io__in_rready = SimpleBus2AXI4Converter_3_io_out_rready; // @[NutShell.scala 121:14]
  assign plic_io__extra_intrVec = REG_1; // @[NutShell.scala 122:29]
  assign SimpleBus2AXI4Converter_3_clock = clock;
  assign SimpleBus2AXI4Converter_3_reset = reset;
  assign SimpleBus2AXI4Converter_3_io_in_req_valid = mmioXbar_io_out_2_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_resp_ready = mmioXbar_io_out_2_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_out_awready = plic_io__in_awready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_wready = plic_io__in_wready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_bvalid = plic_io__in_bvalid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_arready = plic_io__in_arready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_rvalid = plic_io__in_rvalid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_rdata = plic_io__in_rdata; // @[NutShell.scala 121:14]
  always @(posedge clock) begin
    REG <= io_meip; // @[NutShell.scala 122:47]
    REG_1 <= REG; // @[NutShell.scala 122:39]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VGACtrl(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  output        io_in_wready,
  input         io_in_wvalid,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  _T_24 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_25 = io_in_rready & io_in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_25 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_25 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  wire  _T_73 = 4'h0 == io_in_araddr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_74 = 4'h4 == io_in_araddr[3:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_75 = _T_73 ? 32'h190012c : 32'h0; // @[Mux.scala 27:72]
  wire  _T_76 = _T_74 & _T_38; // @[Mux.scala 27:72]
  wire [31:0] _GEN_8 = {{31'd0}, _T_76}; // @[Mux.scala 27:72]
  wire [31:0] _T_77 = _T_75 | _GEN_8; // @[Mux.scala 27:72]
  assign io_in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io_in_wready = io_in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io_in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io_in_arready = io_in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io_in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io_in_rdata = {{32'd0}, _T_77}; // @[RegMap.scala 30:11]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  input  [31:0] io_in_awaddr,
  output        io_in_wready,
  input         io_in_wvalid,
  input  [63:0] io_in_wdata,
  input  [7:0]  io_in_wstrb,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] MEM_0 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_0_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_0_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_0_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_0_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_0_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_0_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_0_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_1 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_1_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_1_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_1_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_1_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_1_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_1_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_1_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_2 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_2_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_2_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_2_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_2_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_2_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_2_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_2_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_3 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_3_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_3_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_3_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_3_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_3_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_3_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_3_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_4 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_4_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_4_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_4_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_4_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_4_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_4_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_4_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_5 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_5_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_5_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_5_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_5_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_5_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_5_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_5_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_6 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_6_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_6_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_6_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_6_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_6_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_6_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_6_MPORT_en; // @[AXI4RAM.scala 63:18]
  reg [7:0] MEM_7 [0:59999]; // @[AXI4RAM.scala 63:18]
  wire  MEM_7_MPORT_1_en; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_7_MPORT_1_addr; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_7_MPORT_1_data; // @[AXI4RAM.scala 63:18]
  wire [7:0] MEM_7_MPORT_data; // @[AXI4RAM.scala 63:18]
  wire [15:0] MEM_7_MPORT_addr; // @[AXI4RAM.scala 63:18]
  wire  MEM_7_MPORT_mask; // @[AXI4RAM.scala 63:18]
  wire  MEM_7_MPORT_en; // @[AXI4RAM.scala 63:18]
  wire  _T_24 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_rvalid ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T_24 | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_36 = REG & (_T_24 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = io_in_rvalid ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _T_36 | _GEN_2; // @[StopWatch.scala 27:{20,24}]
  wire  _T_38 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_39 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _T_38 | _GEN_4; // @[StopWatch.scala 27:{20,24}]
  wire  _T_42 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_39 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _T_42 | _GEN_6; // @[StopWatch.scala 27:{20,24}]
  wire [31:0] _T_45 = io_in_awaddr & 32'h7ffff; // @[AXI4RAM.scala 45:33]
  wire [29:0] _T_47 = {{1'd0}, _T_45[31:3]}; // @[AXI4RAM.scala 48:27]
  wire [28:0] wIdx = _T_47[28:0]; // @[AXI4RAM.scala 48:27]
  wire [31:0] _T_48 = io_in_araddr & 32'h7ffff; // @[AXI4RAM.scala 45:33]
  wire [29:0] _T_50 = {{1'd0}, _T_48[31:3]}; // @[AXI4RAM.scala 49:27]
  wire [28:0] rIdx = _T_50[28:0]; // @[AXI4RAM.scala 49:27]
  wire  _T_52 = wIdx < 29'hea60; // @[AXI4RAM.scala 46:32]
  wire [63:0] rdata = {MEM_7_MPORT_1_data,MEM_6_MPORT_1_data,MEM_5_MPORT_1_data,MEM_4_MPORT_1_data,MEM_3_MPORT_1_data,
    MEM_2_MPORT_1_data,MEM_1_MPORT_1_data,MEM_0_MPORT_1_data}; // @[Cat.scala 30:58]
  reg [63:0] r; // @[Reg.scala 15:16]
  assign MEM_0_MPORT_1_en = 1'h1;
  assign MEM_0_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_0_MPORT_1_data = MEM_0[MEM_0_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_0_MPORT_1_data = MEM_0_MPORT_1_addr >= 16'hea60 ? _RAND_1[7:0] : MEM_0[MEM_0_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_0_MPORT_data = io_in_wdata[7:0];
  assign MEM_0_MPORT_addr = wIdx[15:0];
  assign MEM_0_MPORT_mask = io_in_wstrb[0];
  assign MEM_0_MPORT_en = _T_42 & _T_52;
  assign MEM_1_MPORT_1_en = 1'h1;
  assign MEM_1_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_1_MPORT_1_data = MEM_1[MEM_1_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_1_MPORT_1_data = MEM_1_MPORT_1_addr >= 16'hea60 ? _RAND_3[7:0] : MEM_1[MEM_1_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_1_MPORT_data = io_in_wdata[15:8];
  assign MEM_1_MPORT_addr = wIdx[15:0];
  assign MEM_1_MPORT_mask = io_in_wstrb[1];
  assign MEM_1_MPORT_en = _T_42 & _T_52;
  assign MEM_2_MPORT_1_en = 1'h1;
  assign MEM_2_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_2_MPORT_1_data = MEM_2[MEM_2_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_2_MPORT_1_data = MEM_2_MPORT_1_addr >= 16'hea60 ? _RAND_5[7:0] : MEM_2[MEM_2_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_2_MPORT_data = io_in_wdata[23:16];
  assign MEM_2_MPORT_addr = wIdx[15:0];
  assign MEM_2_MPORT_mask = io_in_wstrb[2];
  assign MEM_2_MPORT_en = _T_42 & _T_52;
  assign MEM_3_MPORT_1_en = 1'h1;
  assign MEM_3_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_3_MPORT_1_data = MEM_3[MEM_3_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_3_MPORT_1_data = MEM_3_MPORT_1_addr >= 16'hea60 ? _RAND_7[7:0] : MEM_3[MEM_3_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_3_MPORT_data = io_in_wdata[31:24];
  assign MEM_3_MPORT_addr = wIdx[15:0];
  assign MEM_3_MPORT_mask = io_in_wstrb[3];
  assign MEM_3_MPORT_en = _T_42 & _T_52;
  assign MEM_4_MPORT_1_en = 1'h1;
  assign MEM_4_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_4_MPORT_1_data = MEM_4[MEM_4_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_4_MPORT_1_data = MEM_4_MPORT_1_addr >= 16'hea60 ? _RAND_9[7:0] : MEM_4[MEM_4_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_4_MPORT_data = io_in_wdata[39:32];
  assign MEM_4_MPORT_addr = wIdx[15:0];
  assign MEM_4_MPORT_mask = io_in_wstrb[4];
  assign MEM_4_MPORT_en = _T_42 & _T_52;
  assign MEM_5_MPORT_1_en = 1'h1;
  assign MEM_5_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_5_MPORT_1_data = MEM_5[MEM_5_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_5_MPORT_1_data = MEM_5_MPORT_1_addr >= 16'hea60 ? _RAND_11[7:0] : MEM_5[MEM_5_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_5_MPORT_data = io_in_wdata[47:40];
  assign MEM_5_MPORT_addr = wIdx[15:0];
  assign MEM_5_MPORT_mask = io_in_wstrb[5];
  assign MEM_5_MPORT_en = _T_42 & _T_52;
  assign MEM_6_MPORT_1_en = 1'h1;
  assign MEM_6_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_6_MPORT_1_data = MEM_6[MEM_6_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_6_MPORT_1_data = MEM_6_MPORT_1_addr >= 16'hea60 ? _RAND_13[7:0] : MEM_6[MEM_6_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_6_MPORT_data = io_in_wdata[55:48];
  assign MEM_6_MPORT_addr = wIdx[15:0];
  assign MEM_6_MPORT_mask = io_in_wstrb[6];
  assign MEM_6_MPORT_en = _T_42 & _T_52;
  assign MEM_7_MPORT_1_en = 1'h1;
  assign MEM_7_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_7_MPORT_1_data = MEM_7[MEM_7_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `else
  assign MEM_7_MPORT_1_data = MEM_7_MPORT_1_addr >= 16'hea60 ? _RAND_15[7:0] : MEM_7[MEM_7_MPORT_1_addr]; // @[AXI4RAM.scala 63:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign MEM_7_MPORT_data = io_in_wdata[63:56];
  assign MEM_7_MPORT_addr = wIdx[15:0];
  assign MEM_7_MPORT_mask = io_in_wstrb[7];
  assign MEM_7_MPORT_en = _T_42 & _T_52;
  assign io_in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io_in_wready = io_in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io_in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io_in_arready = 1'h1; // @[AXI4Slave.scala 71:29]
  assign io_in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io_in_rdata = r; // @[AXI4RAM.scala 71:18]
  always @(posedge clock) begin
    if (MEM_0_MPORT_en & MEM_0_MPORT_mask) begin
      MEM_0[MEM_0_MPORT_addr] <= MEM_0_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_1_MPORT_en & MEM_1_MPORT_mask) begin
      MEM_1[MEM_1_MPORT_addr] <= MEM_1_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_2_MPORT_en & MEM_2_MPORT_mask) begin
      MEM_2[MEM_2_MPORT_addr] <= MEM_2_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_3_MPORT_en & MEM_3_MPORT_mask) begin
      MEM_3[MEM_3_MPORT_addr] <= MEM_3_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_4_MPORT_en & MEM_4_MPORT_mask) begin
      MEM_4[MEM_4_MPORT_addr] <= MEM_4_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_5_MPORT_en & MEM_5_MPORT_mask) begin
      MEM_5[MEM_5_MPORT_addr] <= MEM_5_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_6_MPORT_en & MEM_6_MPORT_mask) begin
      MEM_6[MEM_6_MPORT_addr] <= MEM_6_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (MEM_7_MPORT_en & MEM_7_MPORT_mask) begin
      MEM_7[MEM_7_MPORT_addr] <= MEM_7_MPORT_data; // @[AXI4RAM.scala 63:18]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_24; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    if (REG) begin // @[Reg.scala 16:19]
      r <= rdata; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_3[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_4[initvar] = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_5[initvar] = _RAND_10[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_6[initvar] = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    MEM_7[initvar] = _RAND_14[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_busy = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG_2 = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  r = _RAND_21[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4VGA(
  input         clock,
  input         reset,
  output        io_in_fb_awready,
  input         io_in_fb_awvalid,
  input  [31:0] io_in_fb_awaddr,
  input  [2:0]  io_in_fb_awprot,
  output        io_in_fb_wready,
  input         io_in_fb_wvalid,
  input  [63:0] io_in_fb_wdata,
  input  [7:0]  io_in_fb_wstrb,
  input         io_in_fb_bready,
  output        io_in_fb_bvalid,
  output [1:0]  io_in_fb_bresp,
  output        io_in_fb_arready,
  input         io_in_fb_arvalid,
  input  [31:0] io_in_fb_araddr,
  input  [2:0]  io_in_fb_arprot,
  input         io_in_fb_rready,
  output        io_in_fb_rvalid,
  output [1:0]  io_in_fb_rresp,
  output [63:0] io_in_fb_rdata,
  output        io_in_ctrl_awready,
  input         io_in_ctrl_awvalid,
  input  [31:0] io_in_ctrl_awaddr,
  input  [2:0]  io_in_ctrl_awprot,
  output        io_in_ctrl_wready,
  input         io_in_ctrl_wvalid,
  input  [63:0] io_in_ctrl_wdata,
  input  [7:0]  io_in_ctrl_wstrb,
  input         io_in_ctrl_bready,
  output        io_in_ctrl_bvalid,
  output [1:0]  io_in_ctrl_bresp,
  output        io_in_ctrl_arready,
  input         io_in_ctrl_arvalid,
  input  [31:0] io_in_ctrl_araddr,
  input  [2:0]  io_in_ctrl_arprot,
  input         io_in_ctrl_rready,
  output        io_in_ctrl_rvalid,
  output [1:0]  io_in_ctrl_rresp,
  output [63:0] io_in_ctrl_rdata,
  output [23:0] io_vga_rgb,
  output        io_vga_hsync,
  output        io_vga_vsync,
  output        io_vga_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_clock; // @[AXI4VGA.scala 125:20]
  wire  ctrl_reset; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_awready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_awvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_wready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_wvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_bready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_bvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_arready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_arvalid; // @[AXI4VGA.scala 125:20]
  wire [31:0] ctrl_io_in_araddr; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_rready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_rvalid; // @[AXI4VGA.scala 125:20]
  wire [63:0] ctrl_io_in_rdata; // @[AXI4VGA.scala 125:20]
  wire  fb_clock; // @[AXI4VGA.scala 127:18]
  wire  fb_reset; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_awready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_awvalid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_awaddr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_wready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_wvalid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_wdata; // @[AXI4VGA.scala 127:18]
  wire [7:0] fb_io_in_wstrb; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_bready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_bvalid; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_arready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_arvalid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_araddr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_rready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_rvalid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_rdata; // @[AXI4VGA.scala 127:18]
  wire  _T = io_in_fb_arready & io_in_fb_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_1 = io_in_fb_rready & io_in_fb_rvalid; // @[Decoupled.scala 40:37]
  reg  REG; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_1 ? 1'h0 : REG; // @[StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _T | _GEN_0; // @[StopWatch.scala 27:{20,24}]
  reg [10:0] hCounter; // @[Counter.scala 60:40]
  wire  wrap_wrap = hCounter == 11'h41f; // @[Counter.scala 72:24]
  wire [10:0] _wrap_value_T_1 = hCounter + 11'h1; // @[Counter.scala 76:24]
  reg [9:0] vCounter; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = vCounter == 10'h273; // @[Counter.scala 72:24]
  wire [9:0] _wrap_value_T_3 = vCounter + 10'h1; // @[Counter.scala 76:24]
  wire  hInRange = hCounter >= 11'ha8 & hCounter < 11'h3c8; // @[AXI4VGA.scala 138:63]
  wire  vInRange = vCounter >= 10'h5 & vCounter < 10'h25d; // @[AXI4VGA.scala 138:63]
  wire  hCounterIsOdd = hCounter[0]; // @[AXI4VGA.scala 150:31]
  wire  hCounterIs2 = hCounter[1:0] == 2'h2; // @[AXI4VGA.scala 151:35]
  wire  vCounterIsOdd = vCounter[0]; // @[AXI4VGA.scala 152:31]
  wire  _T_12 = hCounter >= 11'ha7 & hCounter < 11'h3c7; // @[AXI4VGA.scala 138:63]
  wire  nextPixel = _T_12 & vInRange & hCounterIsOdd; // @[AXI4VGA.scala 155:78]
  wire  _T_15 = nextPixel & ~vCounterIsOdd; // @[AXI4VGA.scala 156:41]
  reg [16:0] fbPixelAddrV0; // @[Counter.scala 60:40]
  wire  wrap_wrap_2 = fbPixelAddrV0 == 17'h1d4bf; // @[Counter.scala 72:24]
  wire [16:0] _wrap_value_T_5 = fbPixelAddrV0 + 17'h1; // @[Counter.scala 76:24]
  wire  _T_16 = nextPixel & vCounterIsOdd; // @[AXI4VGA.scala 157:41]
  reg [16:0] fbPixelAddrV1; // @[Counter.scala 60:40]
  wire  wrap_wrap_3 = fbPixelAddrV1 == 17'h1d4bf; // @[Counter.scala 72:24]
  wire [16:0] _wrap_value_T_7 = fbPixelAddrV1 + 17'h1; // @[Counter.scala 76:24]
  wire [16:0] _T_17 = vCounterIsOdd ? fbPixelAddrV1 : fbPixelAddrV0; // @[AXI4VGA.scala 161:35]
  wire [18:0] _T_18 = {_T_17,2'h0}; // @[Cat.scala 30:58]
  reg  REG_1; // @[AXI4VGA.scala 162:31]
  wire  _T_20 = fb_io_in_rready & fb_io_in_rvalid; // @[Decoupled.scala 40:37]
  reg [63:0] r; // @[Reg.scala 27:20]
  wire [63:0] _GEN_14 = _T_20 ? fb_io_in_rdata : r; // @[Reg.scala 28:19 27:20 28:23]
  wire [31:0] color = hCounter[1] ? _GEN_14[63:32] : _GEN_14[31:0]; // @[AXI4VGA.scala 167:23]
  VGACtrl ctrl ( // @[AXI4VGA.scala 125:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_in_awready(ctrl_io_in_awready),
    .io_in_awvalid(ctrl_io_in_awvalid),
    .io_in_wready(ctrl_io_in_wready),
    .io_in_wvalid(ctrl_io_in_wvalid),
    .io_in_bready(ctrl_io_in_bready),
    .io_in_bvalid(ctrl_io_in_bvalid),
    .io_in_arready(ctrl_io_in_arready),
    .io_in_arvalid(ctrl_io_in_arvalid),
    .io_in_araddr(ctrl_io_in_araddr),
    .io_in_rready(ctrl_io_in_rready),
    .io_in_rvalid(ctrl_io_in_rvalid),
    .io_in_rdata(ctrl_io_in_rdata)
  );
  AXI4RAM fb ( // @[AXI4VGA.scala 127:18]
    .clock(fb_clock),
    .reset(fb_reset),
    .io_in_awready(fb_io_in_awready),
    .io_in_awvalid(fb_io_in_awvalid),
    .io_in_awaddr(fb_io_in_awaddr),
    .io_in_wready(fb_io_in_wready),
    .io_in_wvalid(fb_io_in_wvalid),
    .io_in_wdata(fb_io_in_wdata),
    .io_in_wstrb(fb_io_in_wstrb),
    .io_in_bready(fb_io_in_bready),
    .io_in_bvalid(fb_io_in_bvalid),
    .io_in_arready(fb_io_in_arready),
    .io_in_arvalid(fb_io_in_arvalid),
    .io_in_araddr(fb_io_in_araddr),
    .io_in_rready(fb_io_in_rready),
    .io_in_rvalid(fb_io_in_rvalid),
    .io_in_rdata(fb_io_in_rdata)
  );
  assign io_in_fb_awready = fb_io_in_awready; // @[AXI4VGA.scala 130:15]
  assign io_in_fb_wready = fb_io_in_wready; // @[AXI4VGA.scala 131:14]
  assign io_in_fb_bvalid = fb_io_in_bvalid; // @[AXI4VGA.scala 132:14]
  assign io_in_fb_bresp = 2'h0; // @[AXI4VGA.scala 132:14]
  assign io_in_fb_arready = 1'h1; // @[AXI4VGA.scala 133:21]
  assign io_in_fb_rvalid = REG; // @[AXI4VGA.scala 136:20]
  assign io_in_fb_rresp = 2'h0; // @[AXI4VGA.scala 135:24]
  assign io_in_fb_rdata = 64'h0; // @[AXI4VGA.scala 134:24]
  assign io_in_ctrl_awready = ctrl_io_in_awready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_wready = ctrl_io_in_wready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_bvalid = ctrl_io_in_bvalid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_bresp = 2'h0; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_arready = ctrl_io_in_arready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rvalid = ctrl_io_in_rvalid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rresp = 2'h0; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rdata = ctrl_io_in_rdata; // @[AXI4VGA.scala 126:14]
  assign io_vga_rgb = io_vga_valid ? color[23:0] : 24'h0; // @[AXI4VGA.scala 168:20]
  assign io_vga_hsync = hCounter >= 11'h28; // @[AXI4VGA.scala 143:28]
  assign io_vga_vsync = vCounter >= 10'h1; // @[AXI4VGA.scala 144:28]
  assign io_vga_valid = hInRange & vInRange; // @[AXI4VGA.scala 148:28]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_in_awvalid = io_in_ctrl_awvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_wvalid = io_in_ctrl_wvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_bready = io_in_ctrl_bready; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_arvalid = io_in_ctrl_arvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_araddr = io_in_ctrl_araddr; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_rready = io_in_ctrl_rready; // @[AXI4VGA.scala 126:14]
  assign fb_clock = clock;
  assign fb_reset = reset;
  assign fb_io_in_awvalid = io_in_fb_awvalid; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_awaddr = io_in_fb_awaddr; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_wvalid = io_in_fb_wvalid; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_wdata = io_in_fb_wdata; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_wstrb = io_in_fb_wstrb; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_bready = io_in_fb_bready; // @[AXI4VGA.scala 132:14]
  assign fb_io_in_arvalid = REG_1 & hCounterIs2; // @[AXI4VGA.scala 162:43]
  assign fb_io_in_araddr = {{13'd0}, _T_18}; // @[AXI4VGA.scala 161:25]
  assign fb_io_in_rready = 1'h1; // @[AXI4VGA.scala 164:20]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      REG <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG <= _GEN_1;
    end
    if (reset) begin // @[Counter.scala 60:40]
      hCounter <= 11'h0; // @[Counter.scala 60:40]
    end else if (wrap_wrap) begin // @[Counter.scala 86:20]
      hCounter <= 11'h0; // @[Counter.scala 86:28]
    end else begin
      hCounter <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      vCounter <= 10'h0; // @[Counter.scala 60:40]
    end else if (wrap_wrap) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        vCounter <= 10'h0; // @[Counter.scala 86:28]
      end else begin
        vCounter <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      fbPixelAddrV0 <= 17'h0; // @[Counter.scala 60:40]
    end else if (_T_15) begin // @[Counter.scala 118:17]
      if (wrap_wrap_2) begin // @[Counter.scala 86:20]
        fbPixelAddrV0 <= 17'h0; // @[Counter.scala 86:28]
      end else begin
        fbPixelAddrV0 <= _wrap_value_T_5; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      fbPixelAddrV1 <= 17'h0; // @[Counter.scala 60:40]
    end else if (_T_16) begin // @[Counter.scala 118:17]
      if (wrap_wrap_3) begin // @[Counter.scala 86:20]
        fbPixelAddrV1 <= 17'h0; // @[Counter.scala 86:28]
      end else begin
        fbPixelAddrV1 <= _wrap_value_T_7; // @[Counter.scala 76:15]
      end
    end
    REG_1 <= _T_12 & vInRange & hCounterIsOdd; // @[AXI4VGA.scala 155:78]
    if (reset) begin // @[Reg.scala 27:20]
      r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_20) begin // @[Reg.scala 28:19]
      r <= fb_io_in_rdata; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hCounter = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  vCounter = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  fbPixelAddrV0 = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  fbPixelAddrV1 = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  r = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input   clock,
  input   reset
);
  wire  nutshell_clock; // @[TopMain.scala 29:24]
  wire  nutshell_reset; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mem_awaddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_awprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awuser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mem_awlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_awsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_awburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_awlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_awcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_awqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_wready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_wvalid; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mem_wdata; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mem_wstrb; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_wlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_bready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_bvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_bresp; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_bid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_buser; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mem_araddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_arprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_aruser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mem_arlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mem_arsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_arburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_arlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_arcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mem_arqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mem_rresp; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mem_rdata; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_rid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mem_ruser; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mmio_awaddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_awprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awuser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mmio_awlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_awsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_awburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_awlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_awcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_awqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_wready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_wvalid; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mmio_wdata; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mmio_wstrb; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_wlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_bready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_bvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_bresp; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_bid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_buser; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_mmio_araddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_arprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_aruser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_mmio_arlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_mmio_arsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_arburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_arlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_arcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_mmio_arqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rready; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_mmio_rresp; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_mmio_rdata; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_rid; // @[TopMain.scala 29:24]
  wire  nutshell_io_mmio_ruser; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_frontend_awaddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_awprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awuser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_frontend_awlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_awsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_awburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_awlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_awcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_awqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_wready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_wvalid; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_frontend_wdata; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_frontend_wstrb; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_wlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_bready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_bvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_bresp; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_bid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_buser; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arvalid; // @[TopMain.scala 29:24]
  wire [31:0] nutshell_io_frontend_araddr; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_arprot; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_aruser; // @[TopMain.scala 29:24]
  wire [7:0] nutshell_io_frontend_arlen; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_frontend_arsize; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_arburst; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_arlock; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_arcache; // @[TopMain.scala 29:24]
  wire [3:0] nutshell_io_frontend_arqos; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rready; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rvalid; // @[TopMain.scala 29:24]
  wire [1:0] nutshell_io_frontend_rresp; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_frontend_rdata; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rlast; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_rid; // @[TopMain.scala 29:24]
  wire  nutshell_io_frontend_ruser; // @[TopMain.scala 29:24]
  wire [2:0] nutshell_io_meip; // @[TopMain.scala 29:24]
  wire [38:0] nutshell_io_ila_WBUpc; // @[TopMain.scala 29:24]
  wire  nutshell_io_ila_WBUvalid; // @[TopMain.scala 29:24]
  wire  nutshell_io_ila_WBUrfWen; // @[TopMain.scala 29:24]
  wire [4:0] nutshell_io_ila_WBUrfDest; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_ila_WBUrfData; // @[TopMain.scala 29:24]
  wire [63:0] nutshell_io_ila_InstrCnt; // @[TopMain.scala 29:24]
  wire  vga_clock; // @[TopMain.scala 30:19]
  wire  vga_reset; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_awready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_awvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_fb_awaddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_fb_awprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_wready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_wvalid; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_fb_wdata; // @[TopMain.scala 30:19]
  wire [7:0] vga_io_in_fb_wstrb; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_bready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_bvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_fb_bresp; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_arready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_arvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_fb_araddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_fb_arprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_rready; // @[TopMain.scala 30:19]
  wire  vga_io_in_fb_rvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_fb_rresp; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_fb_rdata; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_awready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_awvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_ctrl_awaddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_ctrl_awprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_wready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_wvalid; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_ctrl_wdata; // @[TopMain.scala 30:19]
  wire [7:0] vga_io_in_ctrl_wstrb; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_bready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_bvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_ctrl_bresp; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_arready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_arvalid; // @[TopMain.scala 30:19]
  wire [31:0] vga_io_in_ctrl_araddr; // @[TopMain.scala 30:19]
  wire [2:0] vga_io_in_ctrl_arprot; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_rready; // @[TopMain.scala 30:19]
  wire  vga_io_in_ctrl_rvalid; // @[TopMain.scala 30:19]
  wire [1:0] vga_io_in_ctrl_rresp; // @[TopMain.scala 30:19]
  wire [63:0] vga_io_in_ctrl_rdata; // @[TopMain.scala 30:19]
  wire [23:0] vga_io_vga_rgb; // @[TopMain.scala 30:19]
  wire  vga_io_vga_hsync; // @[TopMain.scala 30:19]
  wire  vga_io_vga_vsync; // @[TopMain.scala 30:19]
  wire  vga_io_vga_valid; // @[TopMain.scala 30:19]
  NutShell nutshell ( // @[TopMain.scala 29:24]
    .clock(nutshell_clock),
    .reset(nutshell_reset),
    .io_mem_awready(nutshell_io_mem_awready),
    .io_mem_awvalid(nutshell_io_mem_awvalid),
    .io_mem_awaddr(nutshell_io_mem_awaddr),
    .io_mem_awprot(nutshell_io_mem_awprot),
    .io_mem_awid(nutshell_io_mem_awid),
    .io_mem_awuser(nutshell_io_mem_awuser),
    .io_mem_awlen(nutshell_io_mem_awlen),
    .io_mem_awsize(nutshell_io_mem_awsize),
    .io_mem_awburst(nutshell_io_mem_awburst),
    .io_mem_awlock(nutshell_io_mem_awlock),
    .io_mem_awcache(nutshell_io_mem_awcache),
    .io_mem_awqos(nutshell_io_mem_awqos),
    .io_mem_wready(nutshell_io_mem_wready),
    .io_mem_wvalid(nutshell_io_mem_wvalid),
    .io_mem_wdata(nutshell_io_mem_wdata),
    .io_mem_wstrb(nutshell_io_mem_wstrb),
    .io_mem_wlast(nutshell_io_mem_wlast),
    .io_mem_bready(nutshell_io_mem_bready),
    .io_mem_bvalid(nutshell_io_mem_bvalid),
    .io_mem_bresp(nutshell_io_mem_bresp),
    .io_mem_bid(nutshell_io_mem_bid),
    .io_mem_buser(nutshell_io_mem_buser),
    .io_mem_arready(nutshell_io_mem_arready),
    .io_mem_arvalid(nutshell_io_mem_arvalid),
    .io_mem_araddr(nutshell_io_mem_araddr),
    .io_mem_arprot(nutshell_io_mem_arprot),
    .io_mem_arid(nutshell_io_mem_arid),
    .io_mem_aruser(nutshell_io_mem_aruser),
    .io_mem_arlen(nutshell_io_mem_arlen),
    .io_mem_arsize(nutshell_io_mem_arsize),
    .io_mem_arburst(nutshell_io_mem_arburst),
    .io_mem_arlock(nutshell_io_mem_arlock),
    .io_mem_arcache(nutshell_io_mem_arcache),
    .io_mem_arqos(nutshell_io_mem_arqos),
    .io_mem_rready(nutshell_io_mem_rready),
    .io_mem_rvalid(nutshell_io_mem_rvalid),
    .io_mem_rresp(nutshell_io_mem_rresp),
    .io_mem_rdata(nutshell_io_mem_rdata),
    .io_mem_rlast(nutshell_io_mem_rlast),
    .io_mem_rid(nutshell_io_mem_rid),
    .io_mem_ruser(nutshell_io_mem_ruser),
    .io_mmio_awready(nutshell_io_mmio_awready),
    .io_mmio_awvalid(nutshell_io_mmio_awvalid),
    .io_mmio_awaddr(nutshell_io_mmio_awaddr),
    .io_mmio_awprot(nutshell_io_mmio_awprot),
    .io_mmio_awid(nutshell_io_mmio_awid),
    .io_mmio_awuser(nutshell_io_mmio_awuser),
    .io_mmio_awlen(nutshell_io_mmio_awlen),
    .io_mmio_awsize(nutshell_io_mmio_awsize),
    .io_mmio_awburst(nutshell_io_mmio_awburst),
    .io_mmio_awlock(nutshell_io_mmio_awlock),
    .io_mmio_awcache(nutshell_io_mmio_awcache),
    .io_mmio_awqos(nutshell_io_mmio_awqos),
    .io_mmio_wready(nutshell_io_mmio_wready),
    .io_mmio_wvalid(nutshell_io_mmio_wvalid),
    .io_mmio_wdata(nutshell_io_mmio_wdata),
    .io_mmio_wstrb(nutshell_io_mmio_wstrb),
    .io_mmio_wlast(nutshell_io_mmio_wlast),
    .io_mmio_bready(nutshell_io_mmio_bready),
    .io_mmio_bvalid(nutshell_io_mmio_bvalid),
    .io_mmio_bresp(nutshell_io_mmio_bresp),
    .io_mmio_bid(nutshell_io_mmio_bid),
    .io_mmio_buser(nutshell_io_mmio_buser),
    .io_mmio_arready(nutshell_io_mmio_arready),
    .io_mmio_arvalid(nutshell_io_mmio_arvalid),
    .io_mmio_araddr(nutshell_io_mmio_araddr),
    .io_mmio_arprot(nutshell_io_mmio_arprot),
    .io_mmio_arid(nutshell_io_mmio_arid),
    .io_mmio_aruser(nutshell_io_mmio_aruser),
    .io_mmio_arlen(nutshell_io_mmio_arlen),
    .io_mmio_arsize(nutshell_io_mmio_arsize),
    .io_mmio_arburst(nutshell_io_mmio_arburst),
    .io_mmio_arlock(nutshell_io_mmio_arlock),
    .io_mmio_arcache(nutshell_io_mmio_arcache),
    .io_mmio_arqos(nutshell_io_mmio_arqos),
    .io_mmio_rready(nutshell_io_mmio_rready),
    .io_mmio_rvalid(nutshell_io_mmio_rvalid),
    .io_mmio_rresp(nutshell_io_mmio_rresp),
    .io_mmio_rdata(nutshell_io_mmio_rdata),
    .io_mmio_rlast(nutshell_io_mmio_rlast),
    .io_mmio_rid(nutshell_io_mmio_rid),
    .io_mmio_ruser(nutshell_io_mmio_ruser),
    .io_frontend_awready(nutshell_io_frontend_awready),
    .io_frontend_awvalid(nutshell_io_frontend_awvalid),
    .io_frontend_awaddr(nutshell_io_frontend_awaddr),
    .io_frontend_awprot(nutshell_io_frontend_awprot),
    .io_frontend_awid(nutshell_io_frontend_awid),
    .io_frontend_awuser(nutshell_io_frontend_awuser),
    .io_frontend_awlen(nutshell_io_frontend_awlen),
    .io_frontend_awsize(nutshell_io_frontend_awsize),
    .io_frontend_awburst(nutshell_io_frontend_awburst),
    .io_frontend_awlock(nutshell_io_frontend_awlock),
    .io_frontend_awcache(nutshell_io_frontend_awcache),
    .io_frontend_awqos(nutshell_io_frontend_awqos),
    .io_frontend_wready(nutshell_io_frontend_wready),
    .io_frontend_wvalid(nutshell_io_frontend_wvalid),
    .io_frontend_wdata(nutshell_io_frontend_wdata),
    .io_frontend_wstrb(nutshell_io_frontend_wstrb),
    .io_frontend_wlast(nutshell_io_frontend_wlast),
    .io_frontend_bready(nutshell_io_frontend_bready),
    .io_frontend_bvalid(nutshell_io_frontend_bvalid),
    .io_frontend_bresp(nutshell_io_frontend_bresp),
    .io_frontend_bid(nutshell_io_frontend_bid),
    .io_frontend_buser(nutshell_io_frontend_buser),
    .io_frontend_arready(nutshell_io_frontend_arready),
    .io_frontend_arvalid(nutshell_io_frontend_arvalid),
    .io_frontend_araddr(nutshell_io_frontend_araddr),
    .io_frontend_arprot(nutshell_io_frontend_arprot),
    .io_frontend_arid(nutshell_io_frontend_arid),
    .io_frontend_aruser(nutshell_io_frontend_aruser),
    .io_frontend_arlen(nutshell_io_frontend_arlen),
    .io_frontend_arsize(nutshell_io_frontend_arsize),
    .io_frontend_arburst(nutshell_io_frontend_arburst),
    .io_frontend_arlock(nutshell_io_frontend_arlock),
    .io_frontend_arcache(nutshell_io_frontend_arcache),
    .io_frontend_arqos(nutshell_io_frontend_arqos),
    .io_frontend_rready(nutshell_io_frontend_rready),
    .io_frontend_rvalid(nutshell_io_frontend_rvalid),
    .io_frontend_rresp(nutshell_io_frontend_rresp),
    .io_frontend_rdata(nutshell_io_frontend_rdata),
    .io_frontend_rlast(nutshell_io_frontend_rlast),
    .io_frontend_rid(nutshell_io_frontend_rid),
    .io_frontend_ruser(nutshell_io_frontend_ruser),
    .io_meip(nutshell_io_meip),
    .io_ila_WBUpc(nutshell_io_ila_WBUpc),
    .io_ila_WBUvalid(nutshell_io_ila_WBUvalid),
    .io_ila_WBUrfWen(nutshell_io_ila_WBUrfWen),
    .io_ila_WBUrfDest(nutshell_io_ila_WBUrfDest),
    .io_ila_WBUrfData(nutshell_io_ila_WBUrfData),
    .io_ila_InstrCnt(nutshell_io_ila_InstrCnt)
  );
  AXI4VGA vga ( // @[TopMain.scala 30:19]
    .clock(vga_clock),
    .reset(vga_reset),
    .io_in_fb_awready(vga_io_in_fb_awready),
    .io_in_fb_awvalid(vga_io_in_fb_awvalid),
    .io_in_fb_awaddr(vga_io_in_fb_awaddr),
    .io_in_fb_awprot(vga_io_in_fb_awprot),
    .io_in_fb_wready(vga_io_in_fb_wready),
    .io_in_fb_wvalid(vga_io_in_fb_wvalid),
    .io_in_fb_wdata(vga_io_in_fb_wdata),
    .io_in_fb_wstrb(vga_io_in_fb_wstrb),
    .io_in_fb_bready(vga_io_in_fb_bready),
    .io_in_fb_bvalid(vga_io_in_fb_bvalid),
    .io_in_fb_bresp(vga_io_in_fb_bresp),
    .io_in_fb_arready(vga_io_in_fb_arready),
    .io_in_fb_arvalid(vga_io_in_fb_arvalid),
    .io_in_fb_araddr(vga_io_in_fb_araddr),
    .io_in_fb_arprot(vga_io_in_fb_arprot),
    .io_in_fb_rready(vga_io_in_fb_rready),
    .io_in_fb_rvalid(vga_io_in_fb_rvalid),
    .io_in_fb_rresp(vga_io_in_fb_rresp),
    .io_in_fb_rdata(vga_io_in_fb_rdata),
    .io_in_ctrl_awready(vga_io_in_ctrl_awready),
    .io_in_ctrl_awvalid(vga_io_in_ctrl_awvalid),
    .io_in_ctrl_awaddr(vga_io_in_ctrl_awaddr),
    .io_in_ctrl_awprot(vga_io_in_ctrl_awprot),
    .io_in_ctrl_wready(vga_io_in_ctrl_wready),
    .io_in_ctrl_wvalid(vga_io_in_ctrl_wvalid),
    .io_in_ctrl_wdata(vga_io_in_ctrl_wdata),
    .io_in_ctrl_wstrb(vga_io_in_ctrl_wstrb),
    .io_in_ctrl_bready(vga_io_in_ctrl_bready),
    .io_in_ctrl_bvalid(vga_io_in_ctrl_bvalid),
    .io_in_ctrl_bresp(vga_io_in_ctrl_bresp),
    .io_in_ctrl_arready(vga_io_in_ctrl_arready),
    .io_in_ctrl_arvalid(vga_io_in_ctrl_arvalid),
    .io_in_ctrl_araddr(vga_io_in_ctrl_araddr),
    .io_in_ctrl_arprot(vga_io_in_ctrl_arprot),
    .io_in_ctrl_rready(vga_io_in_ctrl_rready),
    .io_in_ctrl_rvalid(vga_io_in_ctrl_rvalid),
    .io_in_ctrl_rresp(vga_io_in_ctrl_rresp),
    .io_in_ctrl_rdata(vga_io_in_ctrl_rdata),
    .io_vga_rgb(vga_io_vga_rgb),
    .io_vga_hsync(vga_io_vga_hsync),
    .io_vga_vsync(vga_io_vga_vsync),
    .io_vga_valid(vga_io_vga_valid)
  );
  assign nutshell_clock = clock;
  assign nutshell_reset = reset;
  assign nutshell_io_mem_awready = 1'h0;
  assign nutshell_io_mem_wready = 1'h0;
  assign nutshell_io_mem_bvalid = 1'h0;
  assign nutshell_io_mem_bresp = 2'h0;
  assign nutshell_io_mem_bid = 1'h0;
  assign nutshell_io_mem_buser = 1'h0;
  assign nutshell_io_mem_arready = 1'h0;
  assign nutshell_io_mem_rvalid = 1'h0;
  assign nutshell_io_mem_rresp = 2'h0;
  assign nutshell_io_mem_rdata = 64'h0;
  assign nutshell_io_mem_rlast = 1'h0;
  assign nutshell_io_mem_rid = 1'h0;
  assign nutshell_io_mem_ruser = 1'h0;
  assign nutshell_io_mmio_awready = 1'h0;
  assign nutshell_io_mmio_wready = 1'h0;
  assign nutshell_io_mmio_bvalid = 1'h0;
  assign nutshell_io_mmio_bresp = 2'h0;
  assign nutshell_io_mmio_bid = 1'h0;
  assign nutshell_io_mmio_buser = 1'h0;
  assign nutshell_io_mmio_arready = 1'h0;
  assign nutshell_io_mmio_rvalid = 1'h0;
  assign nutshell_io_mmio_rresp = 2'h0;
  assign nutshell_io_mmio_rdata = 64'h0;
  assign nutshell_io_mmio_rlast = 1'h0;
  assign nutshell_io_mmio_rid = 1'h0;
  assign nutshell_io_mmio_ruser = 1'h0;
  assign nutshell_io_frontend_awvalid = 1'h0;
  assign nutshell_io_frontend_awaddr = 32'h0;
  assign nutshell_io_frontend_awprot = 3'h0;
  assign nutshell_io_frontend_awid = 1'h0;
  assign nutshell_io_frontend_awuser = 1'h0;
  assign nutshell_io_frontend_awlen = 8'h0;
  assign nutshell_io_frontend_awsize = 3'h0;
  assign nutshell_io_frontend_awburst = 2'h0;
  assign nutshell_io_frontend_awlock = 1'h0;
  assign nutshell_io_frontend_awcache = 4'h0;
  assign nutshell_io_frontend_awqos = 4'h0;
  assign nutshell_io_frontend_wvalid = 1'h0;
  assign nutshell_io_frontend_wdata = 64'h0;
  assign nutshell_io_frontend_wstrb = 8'h0;
  assign nutshell_io_frontend_wlast = 1'h0;
  assign nutshell_io_frontend_bready = 1'h0;
  assign nutshell_io_frontend_arvalid = 1'h0;
  assign nutshell_io_frontend_araddr = 32'h0;
  assign nutshell_io_frontend_arprot = 3'h0;
  assign nutshell_io_frontend_arid = 1'h0;
  assign nutshell_io_frontend_aruser = 1'h0;
  assign nutshell_io_frontend_arlen = 8'h0;
  assign nutshell_io_frontend_arsize = 3'h0;
  assign nutshell_io_frontend_arburst = 2'h0;
  assign nutshell_io_frontend_arlock = 1'h0;
  assign nutshell_io_frontend_arcache = 4'h0;
  assign nutshell_io_frontend_arqos = 4'h0;
  assign nutshell_io_frontend_rready = 1'h0;
  assign nutshell_io_meip = 3'h0;
  assign vga_clock = clock;
  assign vga_reset = reset;
  assign vga_io_in_fb_awvalid = 1'h0;
  assign vga_io_in_fb_awaddr = 32'h0;
  assign vga_io_in_fb_awprot = 3'h0;
  assign vga_io_in_fb_wvalid = 1'h0;
  assign vga_io_in_fb_wdata = 64'h0;
  assign vga_io_in_fb_wstrb = 8'h0;
  assign vga_io_in_fb_bready = 1'h0;
  assign vga_io_in_fb_arvalid = 1'h0;
  assign vga_io_in_fb_araddr = 32'h0;
  assign vga_io_in_fb_arprot = 3'h0;
  assign vga_io_in_fb_rready = 1'h0;
  assign vga_io_in_ctrl_awvalid = 1'h0;
  assign vga_io_in_ctrl_awaddr = 32'h0;
  assign vga_io_in_ctrl_awprot = 3'h0;
  assign vga_io_in_ctrl_wvalid = 1'h0;
  assign vga_io_in_ctrl_wdata = 64'h0;
  assign vga_io_in_ctrl_wstrb = 8'h0;
  assign vga_io_in_ctrl_bready = 1'h0;
  assign vga_io_in_ctrl_arvalid = 1'h0;
  assign vga_io_in_ctrl_araddr = 32'h0;
  assign vga_io_in_ctrl_arprot = 3'h0;
  assign vga_io_in_ctrl_rready = 1'h0;
endmodule
module array(
  input  [8:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [72:0] RW0_wdata_0,
  output [72:0] RW0_rdata_0
);
  wire [8:0] array_ext_RW0_addr;
  wire  array_ext_RW0_en;
  wire  array_ext_RW0_clk;
  wire  array_ext_RW0_wmode;
  wire [72:0] array_ext_RW0_wdata;
  wire [72:0] array_ext_RW0_rdata;
  array_ext array_ext (
    .RW0_addr(array_ext_RW0_addr),
    .RW0_en(array_ext_RW0_en),
    .RW0_clk(array_ext_RW0_clk),
    .RW0_wmode(array_ext_RW0_wmode),
    .RW0_wdata(array_ext_RW0_wdata),
    .RW0_rdata(array_ext_RW0_rdata)
  );
  assign array_ext_RW0_clk = RW0_clk;
  assign array_ext_RW0_en = RW0_en;
  assign array_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_ext_RW0_rdata;
  assign array_ext_RW0_wmode = RW0_wmode;
  assign array_ext_RW0_wdata = RW0_wdata_0;
endmodule
module array_0(
  input  [6:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [20:0] RW0_wdata_0,
  input  [20:0] RW0_wdata_1,
  input  [20:0] RW0_wdata_2,
  input  [20:0] RW0_wdata_3,
  output [20:0] RW0_rdata_0,
  output [20:0] RW0_rdata_1,
  output [20:0] RW0_rdata_2,
  output [20:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [6:0] array_0_ext_RW0_addr;
  wire  array_0_ext_RW0_en;
  wire  array_0_ext_RW0_clk;
  wire  array_0_ext_RW0_wmode;
  wire [83:0] array_0_ext_RW0_wdata;
  wire [83:0] array_0_ext_RW0_rdata;
  wire [3:0] array_0_ext_RW0_wmask;
  wire [41:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [41:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_0_ext array_0_ext (
    .RW0_addr(array_0_ext_RW0_addr),
    .RW0_en(array_0_ext_RW0_en),
    .RW0_clk(array_0_ext_RW0_clk),
    .RW0_wmode(array_0_ext_RW0_wmode),
    .RW0_wdata(array_0_ext_RW0_wdata),
    .RW0_rdata(array_0_ext_RW0_rdata),
    .RW0_wmask(array_0_ext_RW0_wmask)
  );
  assign array_0_ext_RW0_clk = RW0_clk;
  assign array_0_ext_RW0_en = RW0_en;
  assign array_0_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_0_ext_RW0_rdata[20:0];
  assign RW0_rdata_1 = array_0_ext_RW0_rdata[41:21];
  assign RW0_rdata_2 = array_0_ext_RW0_rdata[62:42];
  assign RW0_rdata_3 = array_0_ext_RW0_rdata[83:63];
  assign array_0_ext_RW0_wmode = RW0_wmode;
  assign array_0_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_0_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_1(
  input  [9:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [63:0] RW0_wdata_0,
  input  [63:0] RW0_wdata_1,
  input  [63:0] RW0_wdata_2,
  input  [63:0] RW0_wdata_3,
  output [63:0] RW0_rdata_0,
  output [63:0] RW0_rdata_1,
  output [63:0] RW0_rdata_2,
  output [63:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [9:0] array_1_ext_RW0_addr;
  wire  array_1_ext_RW0_en;
  wire  array_1_ext_RW0_clk;
  wire  array_1_ext_RW0_wmode;
  wire [255:0] array_1_ext_RW0_wdata;
  wire [255:0] array_1_ext_RW0_rdata;
  wire [3:0] array_1_ext_RW0_wmask;
  wire [127:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [127:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_1_ext array_1_ext (
    .RW0_addr(array_1_ext_RW0_addr),
    .RW0_en(array_1_ext_RW0_en),
    .RW0_clk(array_1_ext_RW0_clk),
    .RW0_wmode(array_1_ext_RW0_wmode),
    .RW0_wdata(array_1_ext_RW0_wdata),
    .RW0_rdata(array_1_ext_RW0_rdata),
    .RW0_wmask(array_1_ext_RW0_wmask)
  );
  assign array_1_ext_RW0_clk = RW0_clk;
  assign array_1_ext_RW0_en = RW0_en;
  assign array_1_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_1_ext_RW0_rdata[63:0];
  assign RW0_rdata_1 = array_1_ext_RW0_rdata[127:64];
  assign RW0_rdata_2 = array_1_ext_RW0_rdata[191:128];
  assign RW0_rdata_3 = array_1_ext_RW0_rdata[255:192];
  assign array_1_ext_RW0_wmode = RW0_wmode;
  assign array_1_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_1_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_2(
  input  [8:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [18:0] RW0_wdata_0,
  input  [18:0] RW0_wdata_1,
  input  [18:0] RW0_wdata_2,
  input  [18:0] RW0_wdata_3,
  output [18:0] RW0_rdata_0,
  output [18:0] RW0_rdata_1,
  output [18:0] RW0_rdata_2,
  output [18:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [8:0] array_2_ext_RW0_addr;
  wire  array_2_ext_RW0_en;
  wire  array_2_ext_RW0_clk;
  wire  array_2_ext_RW0_wmode;
  wire [75:0] array_2_ext_RW0_wdata;
  wire [75:0] array_2_ext_RW0_rdata;
  wire [3:0] array_2_ext_RW0_wmask;
  wire [37:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [37:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_2_ext array_2_ext (
    .RW0_addr(array_2_ext_RW0_addr),
    .RW0_en(array_2_ext_RW0_en),
    .RW0_clk(array_2_ext_RW0_clk),
    .RW0_wmode(array_2_ext_RW0_wmode),
    .RW0_wdata(array_2_ext_RW0_wdata),
    .RW0_rdata(array_2_ext_RW0_rdata),
    .RW0_wmask(array_2_ext_RW0_wmask)
  );
  assign array_2_ext_RW0_clk = RW0_clk;
  assign array_2_ext_RW0_en = RW0_en;
  assign array_2_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_2_ext_RW0_rdata[18:0];
  assign RW0_rdata_1 = array_2_ext_RW0_rdata[37:19];
  assign RW0_rdata_2 = array_2_ext_RW0_rdata[56:38];
  assign RW0_rdata_3 = array_2_ext_RW0_rdata[75:57];
  assign array_2_ext_RW0_wmode = RW0_wmode;
  assign array_2_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_2_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_3(
  input  [11:0] RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [63:0] RW0_wdata_0,
  input  [63:0] RW0_wdata_1,
  input  [63:0] RW0_wdata_2,
  input  [63:0] RW0_wdata_3,
  output [63:0] RW0_rdata_0,
  output [63:0] RW0_rdata_1,
  output [63:0] RW0_rdata_2,
  output [63:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [11:0] array_3_ext_RW0_addr;
  wire  array_3_ext_RW0_en;
  wire  array_3_ext_RW0_clk;
  wire  array_3_ext_RW0_wmode;
  wire [255:0] array_3_ext_RW0_wdata;
  wire [255:0] array_3_ext_RW0_rdata;
  wire [3:0] array_3_ext_RW0_wmask;
  wire [127:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [127:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_3_ext array_3_ext (
    .RW0_addr(array_3_ext_RW0_addr),
    .RW0_en(array_3_ext_RW0_en),
    .RW0_clk(array_3_ext_RW0_clk),
    .RW0_wmode(array_3_ext_RW0_wmode),
    .RW0_wdata(array_3_ext_RW0_wdata),
    .RW0_rdata(array_3_ext_RW0_rdata),
    .RW0_wmask(array_3_ext_RW0_wmask)
  );
  assign array_3_ext_RW0_clk = RW0_clk;
  assign array_3_ext_RW0_en = RW0_en;
  assign array_3_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_3_ext_RW0_rdata[63:0];
  assign RW0_rdata_1 = array_3_ext_RW0_rdata[127:64];
  assign RW0_rdata_2 = array_3_ext_RW0_rdata[191:128];
  assign RW0_rdata_3 = array_3_ext_RW0_rdata[255:192];
  assign array_3_ext_RW0_wmode = RW0_wmode;
  assign array_3_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_3_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
